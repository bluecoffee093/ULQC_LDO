magic
tech sky130A
magscale 1 2
timestamp 1697794388
<< nmos >>
rect -761 -400 -661 400
rect -603 -400 -503 400
rect -445 -400 -345 400
rect -287 -400 -187 400
rect -129 -400 -29 400
rect 29 -400 129 400
rect 187 -400 287 400
rect 345 -400 445 400
rect 503 -400 603 400
rect 661 -400 761 400
<< ndiff >>
rect -819 388 -761 400
rect -819 -388 -807 388
rect -773 -388 -761 388
rect -819 -400 -761 -388
rect -661 388 -603 400
rect -661 -388 -649 388
rect -615 -388 -603 388
rect -661 -400 -603 -388
rect -503 388 -445 400
rect -503 -388 -491 388
rect -457 -388 -445 388
rect -503 -400 -445 -388
rect -345 388 -287 400
rect -345 -388 -333 388
rect -299 -388 -287 388
rect -345 -400 -287 -388
rect -187 388 -129 400
rect -187 -388 -175 388
rect -141 -388 -129 388
rect -187 -400 -129 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 129 388 187 400
rect 129 -388 141 388
rect 175 -388 187 388
rect 129 -400 187 -388
rect 287 388 345 400
rect 287 -388 299 388
rect 333 -388 345 388
rect 287 -400 345 -388
rect 445 388 503 400
rect 445 -388 457 388
rect 491 -388 503 388
rect 445 -400 503 -388
rect 603 388 661 400
rect 603 -388 615 388
rect 649 -388 661 388
rect 603 -400 661 -388
rect 761 388 819 400
rect 761 -388 773 388
rect 807 -388 819 388
rect 761 -400 819 -388
<< ndiffc >>
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
<< poly >>
rect -761 400 -661 426
rect -603 400 -503 426
rect -445 400 -345 426
rect -287 400 -187 426
rect -129 400 -29 426
rect 29 400 129 426
rect 187 400 287 426
rect 345 400 445 426
rect 503 400 603 426
rect 661 400 761 426
rect -761 -426 -661 -400
rect -603 -426 -503 -400
rect -445 -426 -345 -400
rect -287 -426 -187 -400
rect -129 -426 -29 -400
rect 29 -426 129 -400
rect 187 -426 287 -400
rect 345 -426 445 -400
rect 503 -426 603 -400
rect 661 -426 761 -400
<< locali >>
rect -807 388 -773 404
rect -807 -404 -773 -388
rect -649 388 -615 404
rect -649 -404 -615 -388
rect -491 388 -457 404
rect -491 -404 -457 -388
rect -333 388 -299 404
rect -333 -404 -299 -388
rect -175 388 -141 404
rect -175 -404 -141 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 141 388 175 404
rect 141 -404 175 -388
rect 299 388 333 404
rect 299 -404 333 -388
rect 457 388 491 404
rect 457 -404 491 -388
rect 615 388 649 404
rect 615 -404 649 -388
rect 773 388 807 404
rect 773 -404 807 -388
<< viali >>
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
<< metal1 >>
rect -813 388 -767 400
rect -813 -388 -807 388
rect -773 -388 -767 388
rect -813 -400 -767 -388
rect -655 388 -609 400
rect -655 -388 -649 388
rect -615 -388 -609 388
rect -655 -400 -609 -388
rect -497 388 -451 400
rect -497 -388 -491 388
rect -457 -388 -451 388
rect -497 -400 -451 -388
rect -339 388 -293 400
rect -339 -388 -333 388
rect -299 -388 -293 388
rect -339 -400 -293 -388
rect -181 388 -135 400
rect -181 -388 -175 388
rect -141 -388 -135 388
rect -181 -400 -135 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 135 388 181 400
rect 135 -388 141 388
rect 175 -388 181 388
rect 135 -400 181 -388
rect 293 388 339 400
rect 293 -388 299 388
rect 333 -388 339 388
rect 293 -400 339 -388
rect 451 388 497 400
rect 451 -388 457 388
rect 491 -388 497 388
rect 451 -400 497 -388
rect 609 388 655 400
rect 609 -388 615 388
rect 649 -388 655 388
rect 609 -400 655 -388
rect 767 388 813 400
rect 767 -388 773 388
rect 807 -388 813 388
rect 767 -400 813 -388
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 0.5 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
