* NGSPICE file created from opamp.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_lvt_A3UXRA a_3423_n1000# a_4623_1130# a_1743_1130#
+ a_3135_n1000# a_1503_n3218# a_n3297_1218# a_n4641_1218# a_1215_n3218# a_n1761_1218#
+ a_207_1130# a_n4161_n3218# a_n33_n3218# a_n3921_n1088# a_1119_1218# a_n2289_1022#
+ a_n3345_n1088# a_n3633_1022# a_4239_1130# a_1359_1130# a_3231_n1000# a_n4257_1218#
+ a_2703_1130# a_1311_n3218# a_n1377_1218# a_1023_n3218# a_n2721_1218# a_n465_3240#
+ a_n3249_1022# a_n1713_1022# a_n3153_n1088# a_2319_1130# a_n3969_n1000# a_n2337_1218#
+ a_n1329_1022# a_n4209_1022# a_n3777_n1000# a_n3489_n1000# a_n1857_n3218# a_n1569_n3218#
+ a_n609_n3218# a_n3873_n1000# a_n3585_n1000# a_n1953_n3218# a_n3297_n1000# a_n1665_n3218#
+ a_n1377_n3218# a_n1089_n3218# a_n705_n3218# a_n129_n3218# a_n417_n3218# a_n513_1218#
+ a_n3681_n1000# a_n3393_n1000# a_n1761_n3218# a_n1185_n3218# a_n1473_n3218# a_n753_1130#
+ a_3471_1022# a_n801_n3218# a_n513_n3218# a_4095_1218# a_n129_1218# a_n225_n3218#
+ a_n369_1130# a_3087_1022# a_4431_1022# a_n1281_n3218# a_1551_1022# a_n2385_3240#
+ a_n321_n3218# a_2175_1218# a_4047_1022# a_2799_n1196# a_1167_1022# a_2511_1022#
+ a_n3345_3240# a_3135_1218# a_2127_1022# a_n3393_1218# a_n4305_3240# a_n1425_3240#
+ a_1215_1218# a_2991_n1196# a_63_1218# a_n4353_1218# a_n1473_1218# a_n3729_n1196#
+ a_n4593_1130# a_n1089_1218# a_n2433_1218# a_15_1022# a_n3537_n1196# a_n2673_1130#
+ a_2895_n3306# a_4767_n3218# a_4479_n3218# a_n2049_1218# a_n3921_n1196# a_n4829_1218#
+ a_n2289_1130# a_n3345_n1196# a_n3633_1130# a_n561_1022# a_4575_n3218# a_4287_n3218#
+ a_n3009_1218# a_3183_3240# a_3759_n1088# a_n3249_1130# a_n177_1022# a_n3153_n1196#
+ a_111_3240# a_n1713_1130# a_4671_n3218# a_4383_n3218# a_4095_n3218# a_879_3240#
+ a_n3825_n3306# a_927_n3218# a_4143_3240# a_3567_n1088# a_n3249_n3306# a_639_n3218#
+ a_1263_3240# a_n4209_1130# a_n1329_1130# a_4191_n3218# a_4191_1218# a_n225_1218#
+ a_3951_n1088# a_n3633_n3306# a_735_n3218# a_2223_3240# a_n3057_n3306# a_447_n3218#
+ a_3375_n1088# a_159_n3218# a_2271_1218# a_n3441_n3306# a_831_n3218# a_543_n3218#
+ a_255_n3218# a_3183_n1088# a_3999_n1000# a_3231_1218# a_351_n3218# a_3471_1130#
+ a_3999_1218# a_n4305_n1088# a_927_1218# a_1887_n3218# a_1599_n3218# a_1311_1218#
+ a_n2481_1022# a_3087_1130# a_4431_1130# a_1551_1130# a_n4113_n1088# a_1983_n3218#
+ a_1695_n3218# a_n2097_1022# a_n3441_1022# a_63_n1000# a_4047_1130# a_2511_1130#
+ a_1167_1130# a_n1185_1218# a_n4065_1218# a_n273_3240# a_1791_n3218# a_n3057_1022#
+ a_n4737_n1000# a_n4401_1022# a_n1521_1022# a_n4449_n1000# a_n2817_n3218# a_2127_1130#
+ a_n2529_n3218# a_n2145_1218# a_n4017_1022# a_n1137_1022# a_n4545_n1000# a_n4257_n1000#
+ a_n2913_n3218# a_n2337_n3218# a_n2625_n3218# a_n3105_1218# a_n2049_n3218# a_n1809_n1088#
+ a_n4641_n1000# a_1407_n1000# a_n4353_n1000# a_1119_n1000# a_n2721_n3218# a_n4065_n1000#
+ a_n2433_n3218# a_n2145_n3218# a_15_1130# a_n1617_n1088# a_1503_n1000# a_1215_n1000#
+ a_n4161_n1000# a_n2241_n3218# a_n33_n1000# a_n321_1218# a_n897_n3218# a_n1425_n1088#
+ a_n561_1130# a_1023_n1000# a_1311_n1000# a_3759_n1196# a_975_1022# a_n993_n3218#
+ a_n177_1130# a_n1233_n1088# a_n2193_3240# a_3567_n1196# a_n1041_n1088# a_n3153_3240#
+ a_n1857_n1000# a_3951_n1196# a_n1569_n1000# a_3375_n1196# a_n609_n1000# a_n4113_3240#
+ a_639_1218# a_n1233_3240# a_n1953_n1000# a_n1665_n1000# a_n1377_n1000# a_1023_1218#
+ a_n1089_n1000# a_3183_n1196# a_n705_n1000# a_n417_n1000# a_n1281_1218# a_n4161_1218#
+ a_n129_n1000# a_3855_n3306# a_n1761_n1000# a_3279_n3306# a_n1473_n1000# a_n1185_n1000#
+ a_15_n3306# a_n801_n1000# a_n4305_n1196# a_n513_n1000# a_n225_n1000# a_n2241_1218#
+ a_3663_n3306# a_n2481_1130# a_n1281_n1000# a_3087_n3306# a_4719_n1088# a_n321_n1000#
+ a_n4113_n1196# a_n3201_1218# a_3471_n3306# a_n2097_1130# a_n3969_1218# a_n3441_1130#
+ a_4527_n1088# a_n4209_n3306# a_n3057_1130# a_n4401_1130# a_n1521_1130# a_4335_n1088#
+ a_n4017_n3306# a_687_3240# a_1071_3240# a_n4017_1130# a_n1137_1130# a_n4401_n3306#
+ a_4143_n1088# a_n1809_n1196# a_2031_3240# a_2799_3240# a_n1617_n1196# a_4479_n1000#
+ a_4767_n1000# a_2847_n3218# a_2559_n3218# a_3759_3240# a_n1425_n1196# a_n4689_n1088#
+ a_303_n1088# a_4575_n1000# a_2943_n3218# a_4719_3240# a_4287_n1000# a_2655_n3218#
+ a_1839_3240# a_2367_n3218# a_2079_n3218# a_735_1218# a_1839_n1088# a_n33_1218# a_n1233_n1196#
+ a_n4497_n1088# a_975_1130# a_111_n1088# a_4671_n1000# a_4767_1218# a_4383_n1000#
+ a_2751_n3218# a_1887_1218# a_927_n1000# a_4095_n1000# a_2463_n3218# a_639_n1000#
+ a_n1905_n3306# a_2175_n3218# a_n1329_n3306# a_1647_n1088# a_n1041_n1196# a_4191_n1000#
+ a_2847_1218# a_2271_n3218# a_447_n1000# a_735_n1000# a_n1713_n3306# a_159_n1000#
+ a_1455_n1088# a_n1137_n3306# a_n3009_n3218# a_3807_1218# a_831_n1000# a_543_n1000#
+ a_255_n1000# a_n1521_n3306# a_1263_n1088# a_n3105_n3218# a_n81_n1088# a_351_n1000#
+ a_1071_n1088# a_n3201_n3218# a_n81_3240# a_1599_n1000# a_1887_n1000# a_4719_n1196#
+ a_n849_3240# a_1983_n1000# a_1695_n1000# a_n849_n1088# a_n897_1218# a_4527_n1196#
+ a_1791_n1000# a_n2001_n1088# a_n657_n1088# a_783_1022# a_n2817_n1000# a_n2529_n1000#
+ a_4335_n1196# a_399_1022# a_n2913_n1000# a_n465_n1088# a_n2625_n1000# a_n2337_n1000#
+ a_n2049_n1000# a_4143_n1196# a_831_1218# a_2895_1022# a_n273_n1088# a_n2721_n1000#
+ a_n2433_n1000# a_4239_n3306# a_1983_1218# a_n2145_n1000# a_n1041_3240# a_447_1218#
+ a_3855_1022# a_n4689_3240# a_4623_n3306# a_4479_1218# a_1599_1218# a_4047_n3306#
+ a_2943_1218# a_n2241_n1000# a_n2001_3240# a_n4689_n1196# a_n897_n1000# a_303_n1196#
+ a_1935_1022# a_n2769_3240# a_4431_n3306# a_3903_1218# a_2559_1218# a_1839_n1196#
+ a_n993_n1000# a_n4497_n1196# a_n3729_3240# a_111_n1196# a_3519_1218# a_1647_n1196#
+ a_207_n3306# a_n3777_1218# a_n1809_3240# a_1455_n1196# a_n4829_n3218# a_n4737_1218#
+ a_n1857_1218# a_495_3240# a_n4785_n3306# a_1263_n1196# a_n2817_1218# a_n993_1218#
+ a_2991_3240# a_n81_n1196# a_1935_n3306# a_3807_n3218# a_n4593_n3306# a_1359_n3306#
+ a_3519_n3218# a_1071_n1196# a_879_n1088# a_3951_3240# a_1743_n3306# a_n945_1022#
+ a_3903_n3218# a_3615_n3218# a_1167_n3306# a_3327_n3218# a_3039_n3218# a_3567_3240#
+ a_687_n1088# a_n849_n1196# a_1551_n3306# a_3711_n3218# a_3423_n3218# a_3135_n3218#
+ a_4527_3240# a_2607_n1088# a_1647_3240# a_495_n1088# a_n2001_n1196# a_543_1218#
+ a_n657_n1196# a_783_1130# a_3231_n3218# a_4575_1218# a_1695_1218# a_n609_1218# a_2415_n1088#
+ a_2607_3240# a_159_1218# a_399_1130# a_n465_n1196# a_n3969_n3218# a_2655_1218# a_2223_n1088#
+ a_2895_1130# a_n273_n1196# a_3615_1218# a_n3489_n3218# a_n3777_n3218# a_n4785_1022#
+ a_2031_n1088# a_n945_n3306# a_3855_1130# a_2847_n1000# a_n369_n3306# a_n3873_1218#
+ a_2559_n1000# a_n3873_n3218# a_n2865_1022# a_n3585_n3218# a_n3297_n3218# a_n2769_n1088#
+ a_1935_1130# a_n753_n3306# a_n3489_1218# a_2655_n1000# a_2943_n1000# a_n177_n3306#
+ a_n1953_1218# a_2367_n1000# a_2079_n1000# a_n3681_n3218# a_n3393_n3218# a_n3825_1022#
+ a_n4449_1218# a_n2577_n1088# a_n561_n3306# a_n1569_1218# a_n2913_1218# a_n657_3240#
+ a_2751_n1000# a_2175_n1000# a_2463_n1000# a_n1905_1022# a_n2961_n1088# a_n2529_1218#
+ a_n2385_n1088# a_2271_n1000# a_n3009_n1000# a_591_1022# a_n2193_n1088# a_n3105_n1000#
+ a_n3201_n1000# a_879_n1196# a_4671_1218# a_1791_1218# a_n705_1218# a_255_1218# a_n945_1130#
+ a_3663_1022# a_n4497_3240# a_n2961_3240# a_4287_1218# a_687_n1196# a_2751_1218#
+ a_3279_1022# a_4623_1022# a_1743_1022# a_n2577_3240# a_n3921_3240# a_207_1022# a_2607_n1196#
+ a_2367_1218# a_495_n1196# a_3711_1218# a_4239_1022# a_1359_1022# a_2703_1022# a_n3537_3240#
+ a_2415_n1196# a_3327_1218# a_2319_1022# a_n3585_1218# a_975_n3306# a_n1617_3240#
+ a_399_n3306# a_2223_n1196# a_1407_1218# a_n4545_1218# a_n1665_1218# a_783_n3306#
+ a_2319_n3306# a_n4785_1130# a_2031_n1196# a_2703_n3306# a_n2625_1218# a_591_n3306#
+ a_2127_n3306# a_n2865_1130# a_n2769_n1196# a_3999_n3218# a_2511_n3306# a_n3825_1130#
+ a_n753_1022# a_n2577_n1196# a_3375_3240# a_n369_1022# a_303_3240# a_n1905_1130#
+ a_n2961_n1196# a_n2385_n1196# a_n801_1218# a_4335_3240# a_1455_3240# a_351_1218#
+ a_n4829_n1000# a_2799_n1088# a_63_n3218# a_591_1130# a_n2193_n1196# a_4383_1218#
+ a_n417_1218# a_2415_3240# a_n2865_n3306# a_n4737_n3218# a_n2289_n3306# a_n4449_n3218#
+ a_2463_1218# a_3807_n1000# a_3519_n1000# a_n2673_n3306# a_2991_n1088# a_n4545_n3218#
+ a_n2097_n3306# a_n4257_n3218# a_2079_1218# a_n3729_n1088# a_n4593_1022# a_3423_1218#
+ a_3903_n1000# a_3327_n1000# a_3615_n1000# a_3663_1130# a_3039_n1000# a_1407_n3218#
+ VSUBS a_n2481_n3306# a_n4641_n3218# a_1119_n3218# a_n3681_1218# a_n4065_n3218# a_n4353_n3218#
+ a_3039_1218# a_n3537_n1088# a_1503_1218# a_n2673_1022# a_3711_n1000# a_3279_1130#
X0 a_n321_1218# a_n369_1130# a_n417_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X1 a_2463_n1000# a_2415_n1088# a_2367_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X2 a_n2529_1218# a_n2577_3240# a_n2625_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X3 a_3135_n3218# a_3087_n3306# a_3039_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X4 a_1119_n3218# a_1071_n1196# a_1023_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X5 a_3519_1218# a_3471_1130# a_3423_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X6 a_3135_n1000# a_3087_1022# a_3039_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X7 a_n4641_1218# a_n4689_3240# a_n4737_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X8 a_1503_1218# a_1455_3240# a_1407_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X9 a_n4257_n1000# a_n4305_n1088# a_n4353_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X10 a_1119_n1000# a_1071_n1088# a_1023_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X11 a_n129_n3218# a_n177_n3306# a_n225_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X12 a_543_1218# a_495_3240# a_447_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X13 a_159_n1000# a_111_n1088# a_63_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X14 a_1599_n3218# a_1551_n3306# a_1503_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X15 a_447_n3218# a_399_n3306# a_351_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X16 a_n1185_1218# a_n1233_3240# a_n1281_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X17 a_n2241_n1000# a_n2289_1022# a_n2337_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X18 a_2175_1218# a_2127_1130# a_2079_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X19 a_n3777_n1000# a_n3825_1022# a_n3873_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X20 a_2175_n3218# a_2127_n3306# a_2079_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X21 a_n609_n3218# a_n657_n1196# a_n705_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X22 a_4767_n1000# a_4719_n1088# a_4671_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.1e+12p pd=2.062e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X23 a_n1089_n3218# a_n1137_n3306# a_n1185_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X24 a_n2817_1218# a_n2865_1130# a_n2913_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X25 a_n225_n1000# a_n273_n1088# a_n321_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X26 a_2751_n1000# a_2703_1022# a_2655_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X27 a_4287_n3218# a_4239_n3306# a_4191_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X28 a_3807_1218# a_3759_3240# a_3711_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X29 a_2655_n3218# a_2607_n1196# a_2559_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X30 a_n3489_1218# a_n3537_3240# a_n3585_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X31 a_1791_1218# a_1743_1130# a_1695_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X32 a_1215_n3218# a_1167_n3306# a_1119_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X33 a_831_1218# a_783_1130# a_735_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X34 a_4479_1218# a_4431_1130# a_4383_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X35 a_n4545_n1000# a_n4593_1022# a_n4641_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X36 a_1407_n1000# a_1359_1022# a_1311_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X37 a_4767_n3218# a_4719_n1196# a_4671_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.1e+12p pd=2.062e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X38 a_3231_n3218# a_3183_n1196# a_3135_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X39 a_n1473_1218# a_n1521_1130# a_n1569_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X40 a_447_n1000# a_399_1022# a_351_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X41 a_2463_1218# a_2415_3240# a_2367_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X42 a_n1089_n1000# a_n1137_1022# a_n1185_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X43 a_3327_n3218# a_3279_n3306# a_3231_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X44 a_2079_n1000# a_2031_n1088# a_1983_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X45 a_1695_n3218# a_1647_n1196# a_1599_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X46 a_n225_n3218# a_n273_n1196# a_n321_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X47 a_543_n3218# a_495_n1196# a_447_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X48 a_3135_1218# a_3087_1130# a_3039_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X49 a_n3201_n1000# a_n3249_1022# a_n3297_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X50 a_n4257_1218# a_n4305_3240# a_n4353_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X51 a_1119_1218# a_1071_3240# a_1023_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X52 a_4191_n1000# a_4143_n1088# a_4095_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X53 a_3807_n3218# a_3759_n1196# a_3711_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X54 a_2271_n3218# a_2223_n1196# a_2175_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X55 a_159_1218# a_111_3240# a_63_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X56 a_n513_n1000# a_n561_1022# a_n609_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X57 a_n705_n3218# a_n753_n3306# a_n801_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X58 a_n2241_1218# a_n2289_1130# a_n2337_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X59 a_n1185_n3218# a_n1233_n1196# a_n1281_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X60 a_63_n1000# a_15_1022# a_n33_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X61 a_4383_n3218# a_4335_n1196# a_4287_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X62 a_n3777_1218# a_n3825_1130# a_n3873_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X63 a_1695_n1000# a_1647_n1088# a_1599_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X64 a_2751_n3218# a_2703_n3306# a_2655_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X65 a_4767_1218# a_4719_3240# a_4671_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.1e+12p pd=2.062e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X66 a_735_n1000# a_687_n1088# a_639_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X67 a_n3297_n3218# a_n3345_n1196# a_n3393_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X68 a_n1377_n1000# a_n1425_n1088# a_n1473_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X69 a_n225_1218# a_n273_3240# a_n321_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X70 a_2751_1218# a_2703_1130# a_2655_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X71 a_2367_n1000# a_2319_1022# a_2271_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X72 a_1311_n3218# a_1263_n1196# a_1215_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X73 a_n3777_n3218# a_n3825_n3306# a_n3873_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X74 a_3039_n1000# a_2991_n1088# a_2943_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X75 a_3423_n3218# a_3375_n1196# a_3327_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X76 a_n321_n3218# a_n369_n3306# a_n417_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X77 a_n4545_1218# a_n4593_1130# a_n4641_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X78 a_1407_1218# a_1359_1130# a_1311_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X79 a_n801_n1000# a_n849_n1088# a_n897_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X80 a_1791_n3218# a_1743_n3306# a_1695_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X81 a_n2337_n3218# a_n2385_n1196# a_n2433_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X82 a_447_1218# a_399_1130# a_351_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X83 a_n1089_1218# a_n1137_1130# a_n1185_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X84 a_n2145_n1000# a_n2193_n1088# a_n2241_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X85 a_3999_n1000# a_3951_n1088# a_3903_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X86 a_2079_1218# a_2031_3240# a_1983_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X87 a_n4449_n3218# a_n4497_n1196# a_n4545_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X88 a_3903_n3218# a_3855_n3306# a_3807_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X89 a_n801_n3218# a_n849_n1196# a_n897_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X90 a_1983_n1000# a_1935_1022# a_1887_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X91 a_n1281_n3218# a_n1329_n3306# a_n1377_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X92 a_n2817_n3218# a_n2865_n3306# a_n2913_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X93 a_n3201_1218# a_n3249_1130# a_n3297_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X94 a_4191_1218# a_4143_3240# a_4095_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X95 a_n513_1218# a_n561_1130# a_n609_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X96 a_n129_n1000# a_n177_1022# a_n225_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X97 a_2655_n1000# a_2607_n1088# a_2559_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X98 a_n3393_n3218# a_n3441_n3306# a_n3489_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X99 a_63_1218# a_15_1130# a_n33_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X100 a_1695_1218# a_1647_3240# a_1599_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X101 a_n1761_n1000# a_n1809_n1088# a_n1857_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X102 a_735_1218# a_687_3240# a_639_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X103 a_n4449_n1000# a_n4497_n1088# a_n4545_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X104 a_n1857_n3218# a_n1905_n3306# a_n1953_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X105 a_n3873_n3218# a_n3921_n1196# a_n3969_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X106 a_n1377_1218# a_n1425_3240# a_n1473_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X107 a_2367_1218# a_2319_1130# a_2271_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X108 a_n2433_n1000# a_n2481_1022# a_n2529_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X109 a_n4065_n3218# a_n4113_n1196# a_n4161_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X110 a_3423_n1000# a_3375_n1088# a_3327_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X111 a_n2433_n3218# a_n2481_n3306# a_n2529_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X112 a_n3969_n3218# a_n4017_n3306# a_n4065_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X113 a_3039_1218# a_2991_3240# a_2943_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X114 a_n3105_n1000# a_n3153_n1088# a_n3201_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X115 a_n801_1218# a_n849_3240# a_n897_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X116 a_2943_n1000# a_2895_1022# a_2847_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X117 a_4095_n1000# a_4047_1022# a_3999_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X118 a_n4545_n3218# a_n4593_n3306# a_n4641_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X119 a_n417_n1000# a_n465_n1088# a_n513_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X120 a_n2913_n3218# a_n2961_n1196# a_n3009_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X121 a_n2145_1218# a_n2193_3240# a_n2241_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X122 a_3999_1218# a_3951_3240# a_3903_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X123 a_1983_1218# a_1935_1130# a_1887_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X124 a_n4737_n1000# a_n4785_1022# a_n4829_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.1e+12p ps=2.062e+07u w=1e+07u l=150000u
X125 a_1599_n1000# a_1551_1022# a_1503_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X126 a_n2721_n1000# a_n2769_n1088# a_n2817_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X127 a_639_n1000# a_591_1022# a_543_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X128 a_n129_1218# a_n177_1130# a_n225_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X129 a_2655_1218# a_2607_3240# a_2559_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X130 a_3711_n1000# a_3663_1022# a_3615_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X131 a_n1953_n3218# a_n2001_n1196# a_n2049_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X132 a_n3393_n1000# a_n3441_1022# a_n3489_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X133 a_n4161_n3218# a_n4209_n3306# a_n4257_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X134 a_n1761_1218# a_n1809_3240# a_n1857_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X135 a_4383_n1000# a_4335_n1088# a_4287_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X136 a_n4449_1218# a_n4497_3240# a_n4545_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X137 a_n705_n1000# a_n753_1022# a_n801_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X138 a_159_n3218# a_111_n1196# a_63_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X139 a_n2433_1218# a_n2481_1130# a_n2529_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X140 a_n4641_n3218# a_n4689_n1196# a_n4737_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X141 a_63_n3218# a_15_n3306# a_n33_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X142 a_3423_1218# a_3375_3240# a_3327_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X143 a_n2049_n1000# a_n2097_1022# a_n2145_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X144 a_1887_n1000# a_1839_n1088# a_1791_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X145 a_639_n3218# a_591_n3306# a_543_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X146 a_n3105_1218# a_n3153_3240# a_n3201_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X147 a_2943_1218# a_2895_1130# a_2847_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X148 a_4095_1218# a_4047_1130# a_3999_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X149 a_n4161_n1000# a_n4209_1022# a_n4257_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X150 a_n417_1218# a_n465_3240# a_n513_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X151 a_2559_n1000# a_2511_1022# a_2463_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X152 a_2367_n3218# a_2319_n3306# a_2271_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X153 a_n3681_n1000# a_n3729_n1088# a_n3777_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X154 a_1023_n1000# a_975_1022# a_927_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X155 a_n4737_1218# a_n4785_1130# a_n4829_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.1e+12p ps=2.062e+07u w=1e+07u l=150000u
X156 a_1599_1218# a_1551_1130# a_1503_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X157 a_n1665_n1000# a_n1713_1022# a_n1761_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X158 a_4671_n1000# a_4623_1022# a_4575_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X159 a_4479_n3218# a_4431_n3306# a_4383_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X160 a_2847_n3218# a_2799_n1196# a_2751_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X161 a_n2721_1218# a_n2769_3240# a_n2817_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X162 a_639_1218# a_591_1130# a_543_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X163 a_3711_1218# a_3663_1130# a_3615_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X164 a_n2337_n1000# a_n2385_n1088# a_n2433_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X165 a_3327_n1000# a_3279_1022# a_3231_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X166 a_1407_n3218# a_1359_n3306# a_1311_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X167 a_255_n3218# a_207_n3306# a_159_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X168 a_n3393_1218# a_n3441_1130# a_n3489_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X169 a_4383_1218# a_4335_3240# a_4287_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X170 a_n3009_n1000# a_n3057_1022# a_n3105_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X171 a_1311_n1000# a_1263_n1088# a_1215_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X172 a_n705_1218# a_n753_1130# a_n801_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X173 a_351_n1000# a_303_n1088# a_255_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X174 a_2847_n1000# a_2799_n1088# a_2751_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X175 a_3519_n3218# a_3471_n3306# a_3423_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X176 a_n417_n3218# a_n465_n1196# a_n513_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X177 a_n3969_n1000# a_n4017_1022# a_n4065_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X178 a_n993_n1000# a_n1041_n1088# a_n1089_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X179 a_n33_n1000# a_n81_n1088# a_n129_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X180 a_1887_n3218# a_1839_n1196# a_1791_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X181 a_735_n3218# a_687_n1196# a_639_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X182 a_n2049_1218# a_n2097_1130# a_n2145_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X183 a_n1953_n1000# a_n2001_n1088# a_n2049_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X184 a_4095_n3218# a_4047_n3306# a_3999_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X185 a_1887_1218# a_1839_3240# a_1791_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X186 a_3999_n3218# a_3951_n1196# a_3903_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X187 a_2463_n3218# a_2415_n1196# a_2367_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X188 a_n897_n3218# a_n945_n3306# a_n993_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X189 a_n3009_n3218# a_n3057_n3306# a_n3105_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X190 a_n1377_n3218# a_n1425_n1196# a_n1473_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X191 a_n4161_1218# a_n4209_1130# a_n4257_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X192 a_2559_1218# a_2511_1130# a_2463_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X193 a_n2625_n1000# a_n2673_1022# a_n2721_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X194 a_3615_n1000# a_3567_n1088# a_3519_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X195 a_4575_n3218# a_4527_n1196# a_4479_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X196 a_2943_n3218# a_2895_n3306# a_2847_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X197 a_n3489_n3218# a_n3537_n1196# a_n3585_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X198 a_n3681_1218# a_n3729_3240# a_n3777_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X199 a_1023_1218# a_975_1130# a_927_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X200 a_n1665_1218# a_n1713_1130# a_n1761_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X201 a_4671_1218# a_4623_1130# a_4575_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X202 a_n3297_n1000# a_n3345_n1088# a_n3393_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X203 a_1503_n3218# a_1455_n1196# a_1407_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X204 a_n609_n1000# a_n657_n1088# a_n705_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X205 a_4287_n1000# a_4239_1022# a_4191_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X206 a_351_n3218# a_303_n1196# a_255_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X207 a_n2049_n3218# a_n2097_n3306# a_n2145_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X208 a_n1281_n1000# a_n1329_1022# a_n1377_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X209 a_n2337_1218# a_n2385_3240# a_n2433_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X210 a_2271_n1000# a_2223_n1088# a_2175_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X211 a_3615_n3218# a_3567_n1196# a_3519_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X212 a_3327_1218# a_3279_1130# a_3231_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X213 a_1983_n3218# a_1935_n3306# a_1887_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X214 a_n513_n3218# a_n561_n3306# a_n609_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X215 a_831_n3218# a_783_n3306# a_735_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X216 a_n993_n3218# a_n1041_n1196# a_n1089_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X217 a_n2529_n3218# a_n2577_n1196# a_n2625_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X218 a_n3009_1218# a_n3057_1130# a_n3105_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X219 a_1311_1218# a_1263_3240# a_1215_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X220 a_4191_n3218# a_4143_n1196# a_4095_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X221 a_351_1218# a_303_3240# a_255_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X222 a_2847_1218# a_2799_3240# a_2751_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X223 a_n4065_n1000# a_n4113_n1088# a_n4161_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X224 a_n2913_n1000# a_n2961_n1088# a_n3009_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X225 a_927_n3218# a_879_n1196# a_831_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X226 a_n3969_1218# a_n4017_1130# a_n4065_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X227 a_n993_1218# a_n1041_3240# a_n1089_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X228 a_n33_1218# a_n81_3240# a_n129_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X229 a_3903_n1000# a_3855_1022# a_3807_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X230 a_n3105_n3218# a_n3153_n1196# a_n3201_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X231 a_n1473_n3218# a_n1521_n3306# a_n1569_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X232 a_n1953_1218# a_n2001_3240# a_n2049_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X233 a_n3585_n1000# a_n3633_1022# a_n3681_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X234 a_927_n1000# a_879_n1088# a_831_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X235 a_4671_n3218# a_4623_n3306# a_4575_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X236 a_n1569_n1000# a_n1617_n1088# a_n1665_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X237 a_4575_n1000# a_4527_n1088# a_4479_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X238 a_n1569_n3218# a_n1617_n1196# a_n1665_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X239 a_n897_n1000# a_n945_1022# a_n993_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X240 a_n3585_n3218# a_n3633_n3306# a_n3681_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X241 a_n2625_1218# a_n2673_1130# a_n2721_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X242 a_3615_1218# a_3567_3240# a_3519_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X243 a_n2145_n3218# a_n2193_n1196# a_n2241_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X244 a_3231_n1000# a_3183_n1088# a_3135_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X245 a_n3297_1218# a_n3345_3240# a_n3393_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X246 a_n4353_n1000# a_n4401_1022# a_n4449_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X247 a_1215_n1000# a_1167_1022# a_1119_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X248 a_3711_n3218# a_3663_n3306# a_3615_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X249 a_n4257_n3218# a_n4305_n1196# a_n4353_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X250 a_n609_1218# a_n657_3240# a_n705_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X251 a_4287_1218# a_4239_1130# a_4191_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X252 a_255_n1000# a_207_1022# a_159_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X253 a_n2625_n3218# a_n2673_n3306# a_n2721_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X254 a_n1281_1218# a_n1329_1130# a_n1377_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X255 a_2271_1218# a_2223_3240# a_2175_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X256 a_1023_n3218# a_975_n3306# a_927_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X257 a_n3873_n1000# a_n3921_n1088# a_n3969_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X258 a_n4737_n3218# a_n4785_n3306# a_n4829_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.1e+12p ps=2.062e+07u w=1e+07u l=150000u
X259 a_n3201_n3218# a_n3249_n3306# a_n3297_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X260 a_n1857_n1000# a_n1905_1022# a_n1953_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X261 a_n4065_1218# a_n4113_3240# a_n4161_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X262 a_n2913_1218# a_n2961_3240# a_n3009_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X263 a_n321_n1000# a_n369_1022# a_n417_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X264 a_3903_1218# a_3855_1130# a_3807_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X265 a_n2529_n1000# a_n2577_n1088# a_n2625_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X266 a_n1665_n3218# a_n1713_n3306# a_n1761_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X267 a_n3681_n3218# a_n3729_n1196# a_n3777_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X268 a_3519_n1000# a_3471_1022# a_3423_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X269 a_n3585_1218# a_n3633_1130# a_n3681_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X270 a_927_1218# a_879_3240# a_831_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X271 a_n1569_1218# a_n1617_3240# a_n1665_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X272 a_4575_1218# a_4527_3240# a_4479_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X273 a_n4641_n1000# a_n4689_n1088# a_n4737_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X274 a_1503_n1000# a_1455_n1088# a_1407_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X275 a_n2241_n3218# a_n2289_n3306# a_n2337_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X276 a_n897_1218# a_n945_1130# a_n993_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X277 a_543_n1000# a_495_n1088# a_447_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X278 a_3039_n3218# a_2991_n1196# a_2943_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X279 a_n1185_n1000# a_n1233_n1088# a_n1281_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X280 a_2175_n1000# a_2127_1022# a_2079_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X281 a_n4353_n3218# a_n4401_n3306# a_n4449_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X282 a_n2721_n3218# a_n2769_n1196# a_n2817_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X283 a_3231_1218# a_3183_3240# a_3135_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X284 a_n4353_1218# a_n4401_1130# a_n4449_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X285 a_1215_1218# a_1167_1130# a_1119_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X286 a_255_1218# a_207_1130# a_159_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X287 a_n2817_n1000# a_n2865_1022# a_n2913_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X288 a_2079_n3218# a_2031_n1196# a_1983_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X289 a_3807_n1000# a_3759_n1088# a_3711_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X290 a_n33_n3218# a_n81_n1196# a_n129_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X291 a_n3873_1218# a_n3921_3240# a_n3969_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X292 a_n3489_n1000# a_n3537_n1088# a_n3585_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X293 a_1791_n1000# a_1743_1022# a_1695_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X294 a_n1761_n3218# a_n1809_n1196# a_n1857_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X295 a_n1857_1218# a_n1905_1130# a_n1953_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X296 a_831_n1000# a_783_1022# a_735_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X297 a_4479_n1000# a_4431_1022# a_4383_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X298 a_2559_n3218# a_2511_n3306# a_2463_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X299 a_n1473_n1000# a_n1521_1022# a_n1569_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_477Z4B a_n682_n597# a_n501_n500# a_n855_n500# a_561_n500#
+ a_n383_n500# a_n210_n597# a_n564_n597# a_n737_n500# a_797_n500# a_443_n500# a_380_n597#
+ a_n92_n597# a_n265_n500# a_n446_n597# a_734_n597# a_n619_n500# a_325_n500# a_679_n500#
+ a_n147_n500# a_262_n597# a_n328_n597# a_616_n597# w_n993_n719# a_207_n500# a_144_n597#
+ a_498_n597# a_n29_n500# a_89_n500# a_n800_n597# a_26_n597#
X0 a_325_n500# a_262_n597# a_207_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X1 a_561_n500# a_498_n597# a_443_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X2 a_n265_n500# a_n328_n597# a_n383_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X3 a_797_n500# a_734_n597# a_679_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X4 a_89_n500# a_26_n597# a_n29_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X5 a_207_n500# a_144_n597# a_89_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X6 a_n501_n500# a_n564_n597# a_n619_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X7 a_n147_n500# a_n210_n597# a_n265_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=300000u
X8 a_679_n500# a_616_n597# a_561_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X9 a_n737_n500# a_n800_n597# a_n855_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X10 a_443_n500# a_380_n597# a_325_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X11 a_n383_n500# a_n446_n597# a_n501_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X12 a_n619_n500# a_n682_n597# a_n737_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X13 a_n29_n500# a_n92_n597# a_n147_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
.ends

.subckt sky130_fd_pr__nfet_01v8_Z85A38 a_1261_n500# a_n1319_n500# a_1577_n526# a_n287_n500#
+ a_n1061_n500# a_745_n500# a_29_n526# a_n1777_n526# a_n745_n526# a_1777_n500# a_n2351_n500#
+ a_803_n526# a_n2035_n526# a_229_n500# a_n1577_n500# a_2035_n500# a_1835_n526# a_n229_n526#
+ a_n545_n500# a_287_n526# a_n1003_n526# a_2093_n526# a_1003_n500# a_1319_n526# a_n2293_n526#
+ a_1061_n526# a_n29_n500# a_487_n500# a_2293_n500# a_n1835_n500# a_n1519_n526# a_n487_n526#
+ a_n1261_n526# a_1519_n500# a_n803_n500# a_545_n526# a_n2093_n500# VSUBS
X0 a_n1577_n500# a_n1777_n526# a_n1835_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_1519_n500# a_1319_n526# a_1261_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X2 a_n1061_n500# a_n1261_n526# a_n1319_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_1003_n500# a_803_n526# a_745_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X4 a_487_n500# a_287_n526# a_229_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X5 a_745_n500# a_545_n526# a_487_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X6 a_2035_n500# a_1835_n526# a_1777_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X7 a_1777_n500# a_1577_n526# a_1519_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 a_1261_n500# a_1061_n526# a_1003_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X9 a_n1835_n500# a_n2035_n526# a_n2093_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X10 a_n2093_n500# a_n2293_n526# a_n2351_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X11 a_n29_n500# a_n229_n526# a_n287_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X12 a_229_n500# a_29_n526# a_n29_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X13 a_n1319_n500# a_n1519_n526# a_n1577_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X14 a_n545_n500# a_n745_n526# a_n803_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X15 a_2293_n500# a_2093_n526# a_2035_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X16 a_n803_n500# a_n1003_n526# a_n1061_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X17 a_n287_n500# a_n487_n526# a_n545_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_U3DWQW a_n345_n800# a_129_n800# a_n503_n800# a_29_n826#
+ a_n661_n800# a_n129_n826# a_287_n800# a_187_n826# a_n287_n826# a_445_n800# a_345_n826#
+ a_n445_n826# a_603_n800# a_503_n826# a_n603_n826# a_761_n800# a_661_n826# a_n29_n800#
+ a_n761_n826# a_n187_n800# a_n819_n800# VSUBS
X0 a_n661_n800# a_n761_n826# a_n819_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X1 a_n187_n800# a_n287_n826# a_n345_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X2 a_761_n800# a_661_n826# a_603_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X3 a_287_n800# a_187_n826# a_129_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X4 a_n345_n800# a_n445_n826# a_n503_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X5 a_129_n800# a_29_n826# a_n29_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X6 a_445_n800# a_345_n826# a_287_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=500000u
X7 a_n503_n800# a_n603_n826# a_n661_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X8 a_n29_n800# a_n129_n826# a_n187_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X9 a_603_n800# a_503_n826# a_445_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_2J7QF2 a_147_n526# a_n501_n500# a_561_n500# a_n383_n500#
+ a_29_n526# a_n737_n500# a_n561_n526# a_443_n500# a_n265_n500# a_n443_n526# a_n619_n500#
+ a_325_n500# a_501_n526# a_679_n500# a_n147_n500# a_n325_n526# a_383_n526# a_n679_n526#
+ a_207_n500# a_n29_n500# a_n207_n526# a_265_n526# a_619_n526# a_89_n500# a_n89_n526#
+ VSUBS
X0 a_n383_n500# a_n443_n526# a_n501_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X1 a_n619_n500# a_n679_n526# a_n737_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X2 a_n29_n500# a_n89_n526# a_n147_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X3 a_325_n500# a_265_n526# a_207_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X4 a_n265_n500# a_n325_n526# a_n383_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=300000u
X5 a_561_n500# a_501_n526# a_443_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X6 a_89_n500# a_29_n526# a_n29_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=300000u
X7 a_207_n500# a_147_n526# a_89_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X8 a_n501_n500# a_n561_n526# a_n619_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X9 a_n147_n500# a_n207_n526# a_n265_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X10 a_679_n500# a_619_n526# a_561_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=300000u
X11 a_443_n500# a_383_n526# a_325_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
.ends

.subckt opamp POS NEG VDD VSS BIAS_CUR EA_OUT
Xsky130_fd_pr__nfet_01v8_lvt_A3UXRA_0 VSS VSS VSS P1 VSS VSS VSS P1 VSS VSS P1 VSS
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS P1 VSS
+ VSS VSS P1 VSS P1 VSS VSS VSS P1 VSS VSS P1 VSS P1 P1 P1 VSS P1 VSS P1 VSS VSS P1
+ VSS VSS VSS P1 P1 P1 VSS VSS VSS VSS P1 VSS VSS P1 P1 VSS VSS VSS VSS VSS P1 VSS
+ P1 VSS VSS P1 VSS P1 P1 P1 VSS VSS P1 P1 VSS VSS VSS VSS VSS P1 P1 VSS VSS VSS VSS
+ VSS VSS VSS P1 P1 VSS VSS VSS VSS VSS VSS VSS P1 VSS P1 VSS VSS VSS VSS VSS VSS
+ P1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS P1 VSS P1 VSS
+ VSS VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS P1 VSS
+ VSS VSS VSS VSS VSS P1 VSS P1 VSS VSS VSS P1 VSS VSS VSS VSS VSS P1 VSS VSS VSS
+ P1 VSS P1 VSS VSS P1 P1 VSS VSS VSS P1 VSS VSS VSS VSS P1 P1 P1 VSS P1 P1 VSS VSS
+ P1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS P1 VSS VSS P1
+ VSS P1 P1 VSS P1 VSS P1 P1 P1 VSS VSS VSS P1 VSS VSS VSS VSS P1 VSS P1 VSS VSS P1
+ VSS VSS P1 VSS P1 VSS VSS P1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS
+ VSS VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS VSS VSS VSS P1 VSS P1 VSS VSS P1 VSS VSS
+ VSS VSS VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS P1 VSS P1 VSS P1 VSS VSS VSS VSS VSS
+ VSS P1 VSS VSS VSS VSS VSS P1 VSS P1 VSS P1 VSS VSS VSS VSS VSS VSS P1 VSS P1 VSS
+ VSS VSS P1 VSS VSS P1 VSS P1 VSS VSS VSS P1 VSS VSS VSS VSS VSS P1 VSS P1 VSS P1
+ VSS VSS VSS P1 VSS P1 VSS VSS P1 VSS VSS VSS P1 P1 VSS P1 P1 VSS VSS P1 VSS VSS
+ VSS VSS P1 P1 VSS VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS VSS P1 P1 VSS VSS VSS P1
+ VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS VSS VSS
+ VSS P1 VSS P1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS
+ P1 VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS
+ VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS P1 VSS VSS VSS VSS VSS VSS VSS P1 P1 VSS VSS
+ VSS VSS VSS VSS P1 VSS VSS VSS P1 VSS P1 P1 P1 P1 VSS VSS VSS VSS P1 VSS P1 VSS
+ VSS VSS VSS VSS VSS VSS P1 VSS P1 VSS VSS VSS VSS VSS P1 VSS P1 VSS VSS VSS VSS
+ P1 P1 P1 VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS
+ P1 VSS VSS P1 VSS VSS VSS VSS VSS VSS P1 P1 VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS
+ P1 VSS VSS VSS VSS P1 VSS sky130_fd_pr__nfet_01v8_lvt_A3UXRA
Xsky130_fd_pr__pfet_01v8_477Z4B_0 NEG_D NEG_2 VDD VDD VDD NEG_D NEG_D NEG_D VDD NEG_2
+ NEG_D NEG_D NEG_D NEG_D VDD VDD VDD NEG_D VDD NEG_D NEG_D NEG_D VDD NEG_D NEG_D
+ NEG_D NEG_2 VDD VDD NEG_D sky130_fd_pr__pfet_01v8_477Z4B
Xsky130_fd_pr__pfet_01v8_477Z4B_1 POS_D EA_OUT VDD VDD VDD POS_D POS_D POS_D VDD EA_OUT
+ POS_D POS_D POS_D POS_D VDD VDD VDD POS_D VDD POS_D POS_D POS_D VDD POS_D POS_D
+ POS_D EA_OUT VDD VDD POS_D sky130_fd_pr__pfet_01v8_477Z4B
Xsky130_fd_pr__nfet_01v8_Z85A38_0 VSS VSS BIAS_CUR VSS P1 VSS BIAS_CUR BIAS_CUR BIAS_CUR
+ VSS VSS BIAS_CUR BIAS_CUR VSS BIAS_CUR P1 BIAS_CUR BIAS_CUR BIAS_CUR BIAS_CUR BIAS_CUR
+ VSS P1 BIAS_CUR VSS BIAS_CUR P1 BIAS_CUR VSS VSS BIAS_CUR BIAS_CUR BIAS_CUR BIAS_CUR
+ VSS BIAS_CUR P1 VSS sky130_fd_pr__nfet_01v8_Z85A38
Xsky130_fd_pr__nfet_01v8_U3DWQW_0 POS_D P1 P1 NEG NEG_D NEG POS_D POS POS P1 POS POS
+ NEG_D NEG NEG P1 P1 NEG_D P1 P1 P1 VSS sky130_fd_pr__nfet_01v8_U3DWQW
Xsky130_fd_pr__nfet_01v8_2J7QF2_0 NEG_2 VSS EA_OUT EA_OUT NEG_2 VSS NEG_2 VSS VSS
+ NEG_2 NEG_2 NEG_2 NEG_2 VSS NEG_2 NEG_2 NEG_2 NEG_2 VSS VSS NEG_2 NEG_2 NEG_2 EA_OUT
+ NEG_2 VSS sky130_fd_pr__nfet_01v8_2J7QF2
.ends

