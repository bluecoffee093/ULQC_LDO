magic
tech sky130A
magscale 1 2
timestamp 1697794388
<< error_p >>
rect -442 481 -384 487
rect -324 481 -266 487
rect -206 481 -148 487
rect -88 481 -30 487
rect 30 481 88 487
rect 148 481 206 487
rect 266 481 324 487
rect 384 481 442 487
rect -442 447 -430 481
rect -324 447 -312 481
rect -206 447 -194 481
rect -88 447 -76 481
rect 30 447 42 481
rect 148 447 160 481
rect 266 447 278 481
rect 384 447 396 481
rect -442 441 -384 447
rect -324 441 -266 447
rect -206 441 -148 447
rect -88 441 -30 447
rect 30 441 88 447
rect 148 441 206 447
rect 266 441 324 447
rect 384 441 442 447
rect -442 -447 -384 -441
rect -324 -447 -266 -441
rect -206 -447 -148 -441
rect -88 -447 -30 -441
rect 30 -447 88 -441
rect 148 -447 206 -441
rect 266 -447 324 -441
rect 384 -447 442 -441
rect -442 -481 -430 -447
rect -324 -481 -312 -447
rect -206 -481 -194 -447
rect -88 -481 -76 -447
rect 30 -481 42 -447
rect 148 -481 160 -447
rect 266 -481 278 -447
rect 384 -481 396 -447
rect -442 -487 -384 -481
rect -324 -487 -266 -481
rect -206 -487 -148 -481
rect -88 -487 -30 -481
rect 30 -487 88 -481
rect 148 -487 206 -481
rect 266 -487 324 -481
rect 384 -487 442 -481
<< nwell >>
rect -537 -500 537 500
<< pmos >>
rect -443 -400 -383 400
rect -325 -400 -265 400
rect -207 -400 -147 400
rect -89 -400 -29 400
rect 29 -400 89 400
rect 147 -400 207 400
rect 265 -400 325 400
rect 383 -400 443 400
<< pdiff >>
rect -501 388 -443 400
rect -501 -388 -489 388
rect -455 -388 -443 388
rect -501 -400 -443 -388
rect -383 388 -325 400
rect -383 -388 -371 388
rect -337 -388 -325 388
rect -383 -400 -325 -388
rect -265 388 -207 400
rect -265 -388 -253 388
rect -219 -388 -207 388
rect -265 -400 -207 -388
rect -147 388 -89 400
rect -147 -388 -135 388
rect -101 -388 -89 388
rect -147 -400 -89 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 89 388 147 400
rect 89 -388 101 388
rect 135 -388 147 388
rect 89 -400 147 -388
rect 207 388 265 400
rect 207 -388 219 388
rect 253 -388 265 388
rect 207 -400 265 -388
rect 325 388 383 400
rect 325 -388 337 388
rect 371 -388 383 388
rect 325 -400 383 -388
rect 443 388 501 400
rect 443 -388 455 388
rect 489 -388 501 388
rect 443 -400 501 -388
<< pdiffc >>
rect -489 -388 -455 388
rect -371 -388 -337 388
rect -253 -388 -219 388
rect -135 -388 -101 388
rect -17 -388 17 388
rect 101 -388 135 388
rect 219 -388 253 388
rect 337 -388 371 388
rect 455 -388 489 388
<< poly >>
rect -446 481 -380 497
rect -446 447 -430 481
rect -396 447 -380 481
rect -446 431 -380 447
rect -328 481 -262 497
rect -328 447 -312 481
rect -278 447 -262 481
rect -328 431 -262 447
rect -210 481 -144 497
rect -210 447 -194 481
rect -160 447 -144 481
rect -210 431 -144 447
rect -92 481 -26 497
rect -92 447 -76 481
rect -42 447 -26 481
rect -92 431 -26 447
rect 26 481 92 497
rect 26 447 42 481
rect 76 447 92 481
rect 26 431 92 447
rect 144 481 210 497
rect 144 447 160 481
rect 194 447 210 481
rect 144 431 210 447
rect 262 481 328 497
rect 262 447 278 481
rect 312 447 328 481
rect 262 431 328 447
rect 380 481 446 497
rect 380 447 396 481
rect 430 447 446 481
rect 380 431 446 447
rect -443 400 -383 431
rect -325 400 -265 431
rect -207 400 -147 431
rect -89 400 -29 431
rect 29 400 89 431
rect 147 400 207 431
rect 265 400 325 431
rect 383 400 443 431
rect -443 -431 -383 -400
rect -325 -431 -265 -400
rect -207 -431 -147 -400
rect -89 -431 -29 -400
rect 29 -431 89 -400
rect 147 -431 207 -400
rect 265 -431 325 -400
rect 383 -431 443 -400
rect -446 -447 -380 -431
rect -446 -481 -430 -447
rect -396 -481 -380 -447
rect -446 -497 -380 -481
rect -328 -447 -262 -431
rect -328 -481 -312 -447
rect -278 -481 -262 -447
rect -328 -497 -262 -481
rect -210 -447 -144 -431
rect -210 -481 -194 -447
rect -160 -481 -144 -447
rect -210 -497 -144 -481
rect -92 -447 -26 -431
rect -92 -481 -76 -447
rect -42 -481 -26 -447
rect -92 -497 -26 -481
rect 26 -447 92 -431
rect 26 -481 42 -447
rect 76 -481 92 -447
rect 26 -497 92 -481
rect 144 -447 210 -431
rect 144 -481 160 -447
rect 194 -481 210 -447
rect 144 -497 210 -481
rect 262 -447 328 -431
rect 262 -481 278 -447
rect 312 -481 328 -447
rect 262 -497 328 -481
rect 380 -447 446 -431
rect 380 -481 396 -447
rect 430 -481 446 -447
rect 380 -497 446 -481
<< polycont >>
rect -430 447 -396 481
rect -312 447 -278 481
rect -194 447 -160 481
rect -76 447 -42 481
rect 42 447 76 481
rect 160 447 194 481
rect 278 447 312 481
rect 396 447 430 481
rect -430 -481 -396 -447
rect -312 -481 -278 -447
rect -194 -481 -160 -447
rect -76 -481 -42 -447
rect 42 -481 76 -447
rect 160 -481 194 -447
rect 278 -481 312 -447
rect 396 -481 430 -447
<< locali >>
rect -446 447 -430 481
rect -396 447 -380 481
rect -328 447 -312 481
rect -278 447 -262 481
rect -210 447 -194 481
rect -160 447 -144 481
rect -92 447 -76 481
rect -42 447 -26 481
rect 26 447 42 481
rect 76 447 92 481
rect 144 447 160 481
rect 194 447 210 481
rect 262 447 278 481
rect 312 447 328 481
rect 380 447 396 481
rect 430 447 446 481
rect -489 388 -455 404
rect -489 -404 -455 -388
rect -371 388 -337 404
rect -371 -404 -337 -388
rect -253 388 -219 404
rect -253 -404 -219 -388
rect -135 388 -101 404
rect -135 -404 -101 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 101 388 135 404
rect 101 -404 135 -388
rect 219 388 253 404
rect 219 -404 253 -388
rect 337 388 371 404
rect 337 -404 371 -388
rect 455 388 489 404
rect 455 -404 489 -388
rect -446 -481 -430 -447
rect -396 -481 -380 -447
rect -328 -481 -312 -447
rect -278 -481 -262 -447
rect -210 -481 -194 -447
rect -160 -481 -144 -447
rect -92 -481 -76 -447
rect -42 -481 -26 -447
rect 26 -481 42 -447
rect 76 -481 92 -447
rect 144 -481 160 -447
rect 194 -481 210 -447
rect 262 -481 278 -447
rect 312 -481 328 -447
rect 380 -481 396 -447
rect 430 -481 446 -447
<< viali >>
rect -430 447 -396 481
rect -312 447 -278 481
rect -194 447 -160 481
rect -76 447 -42 481
rect 42 447 76 481
rect 160 447 194 481
rect 278 447 312 481
rect 396 447 430 481
rect -489 -388 -455 388
rect -371 -388 -337 388
rect -253 -388 -219 388
rect -135 -388 -101 388
rect -17 -388 17 388
rect 101 -388 135 388
rect 219 -388 253 388
rect 337 -388 371 388
rect 455 -388 489 388
rect -430 -481 -396 -447
rect -312 -481 -278 -447
rect -194 -481 -160 -447
rect -76 -481 -42 -447
rect 42 -481 76 -447
rect 160 -481 194 -447
rect 278 -481 312 -447
rect 396 -481 430 -447
<< metal1 >>
rect -442 481 -384 487
rect -442 447 -430 481
rect -396 447 -384 481
rect -442 441 -384 447
rect -324 481 -266 487
rect -324 447 -312 481
rect -278 447 -266 481
rect -324 441 -266 447
rect -206 481 -148 487
rect -206 447 -194 481
rect -160 447 -148 481
rect -206 441 -148 447
rect -88 481 -30 487
rect -88 447 -76 481
rect -42 447 -30 481
rect -88 441 -30 447
rect 30 481 88 487
rect 30 447 42 481
rect 76 447 88 481
rect 30 441 88 447
rect 148 481 206 487
rect 148 447 160 481
rect 194 447 206 481
rect 148 441 206 447
rect 266 481 324 487
rect 266 447 278 481
rect 312 447 324 481
rect 266 441 324 447
rect 384 481 442 487
rect 384 447 396 481
rect 430 447 442 481
rect 384 441 442 447
rect -495 388 -449 400
rect -495 -388 -489 388
rect -455 -388 -449 388
rect -495 -400 -449 -388
rect -377 388 -331 400
rect -377 -388 -371 388
rect -337 -388 -331 388
rect -377 -400 -331 -388
rect -259 388 -213 400
rect -259 -388 -253 388
rect -219 -388 -213 388
rect -259 -400 -213 -388
rect -141 388 -95 400
rect -141 -388 -135 388
rect -101 -388 -95 388
rect -141 -400 -95 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 95 388 141 400
rect 95 -388 101 388
rect 135 -388 141 388
rect 95 -400 141 -388
rect 213 388 259 400
rect 213 -388 219 388
rect 253 -388 259 388
rect 213 -400 259 -388
rect 331 388 377 400
rect 331 -388 337 388
rect 371 -388 377 388
rect 331 -400 377 -388
rect 449 388 495 400
rect 449 -388 455 388
rect 489 -388 495 388
rect 449 -400 495 -388
rect -442 -447 -384 -441
rect -442 -481 -430 -447
rect -396 -481 -384 -447
rect -442 -487 -384 -481
rect -324 -447 -266 -441
rect -324 -481 -312 -447
rect -278 -481 -266 -447
rect -324 -487 -266 -481
rect -206 -447 -148 -441
rect -206 -481 -194 -447
rect -160 -481 -148 -447
rect -206 -487 -148 -481
rect -88 -447 -30 -441
rect -88 -481 -76 -447
rect -42 -481 -30 -447
rect -88 -487 -30 -481
rect 30 -447 88 -441
rect 30 -481 42 -447
rect 76 -481 88 -447
rect 30 -487 88 -481
rect 148 -447 206 -441
rect 148 -481 160 -447
rect 194 -481 206 -447
rect 148 -487 206 -481
rect 266 -447 324 -441
rect 266 -481 278 -447
rect 312 -481 324 -447
rect 266 -487 324 -481
rect 384 -447 442 -441
rect 384 -481 396 -447
rect 430 -481 442 -447
rect 384 -487 442 -481
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4 l 0.3 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
