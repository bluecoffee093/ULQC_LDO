magic
tech sky130A
magscale 1 2
timestamp 1697894789
<< nmos >>
rect -761 -800 -661 800
rect -603 -800 -503 800
rect -445 -800 -345 800
rect -287 -800 -187 800
rect -129 -800 -29 800
rect 29 -800 129 800
rect 187 -800 287 800
rect 345 -800 445 800
rect 503 -800 603 800
rect 661 -800 761 800
<< ndiff >>
rect -819 788 -761 800
rect -819 -788 -807 788
rect -773 -788 -761 788
rect -819 -800 -761 -788
rect -661 788 -603 800
rect -661 -788 -649 788
rect -615 -788 -603 788
rect -661 -800 -603 -788
rect -503 788 -445 800
rect -503 -788 -491 788
rect -457 -788 -445 788
rect -503 -800 -445 -788
rect -345 788 -287 800
rect -345 -788 -333 788
rect -299 -788 -287 788
rect -345 -800 -287 -788
rect -187 788 -129 800
rect -187 -788 -175 788
rect -141 -788 -129 788
rect -187 -800 -129 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 129 788 187 800
rect 129 -788 141 788
rect 175 -788 187 788
rect 129 -800 187 -788
rect 287 788 345 800
rect 287 -788 299 788
rect 333 -788 345 788
rect 287 -800 345 -788
rect 445 788 503 800
rect 445 -788 457 788
rect 491 -788 503 788
rect 445 -800 503 -788
rect 603 788 661 800
rect 603 -788 615 788
rect 649 -788 661 788
rect 603 -800 661 -788
rect 761 788 819 800
rect 761 -788 773 788
rect 807 -788 819 788
rect 761 -800 819 -788
<< ndiffc >>
rect -807 -788 -773 788
rect -649 -788 -615 788
rect -491 -788 -457 788
rect -333 -788 -299 788
rect -175 -788 -141 788
rect -17 -788 17 788
rect 141 -788 175 788
rect 299 -788 333 788
rect 457 -788 491 788
rect 615 -788 649 788
rect 773 -788 807 788
<< poly >>
rect -761 800 -661 826
rect -603 800 -503 826
rect -445 800 -345 826
rect -287 800 -187 826
rect -129 800 -29 826
rect 29 800 129 826
rect 187 800 287 826
rect 345 800 445 826
rect 503 800 603 826
rect 661 800 761 826
rect -761 -826 -661 -800
rect -603 -826 -503 -800
rect -445 -826 -345 -800
rect -287 -826 -187 -800
rect -129 -826 -29 -800
rect 29 -826 129 -800
rect 187 -826 287 -800
rect 345 -826 445 -800
rect 503 -826 603 -800
rect 661 -826 761 -800
<< locali >>
rect -807 788 -773 804
rect -807 -804 -773 -788
rect -649 788 -615 804
rect -649 -804 -615 -788
rect -491 788 -457 804
rect -491 -804 -457 -788
rect -333 788 -299 804
rect -333 -804 -299 -788
rect -175 788 -141 804
rect -175 -804 -141 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 141 788 175 804
rect 141 -804 175 -788
rect 299 788 333 804
rect 299 -804 333 -788
rect 457 788 491 804
rect 457 -804 491 -788
rect 615 788 649 804
rect 615 -804 649 -788
rect 773 788 807 804
rect 773 -804 807 -788
<< viali >>
rect -807 -788 -773 788
rect -649 -788 -615 788
rect -491 -788 -457 788
rect -333 -788 -299 788
rect -175 -788 -141 788
rect -17 -788 17 788
rect 141 -788 175 788
rect 299 -788 333 788
rect 457 -788 491 788
rect 615 -788 649 788
rect 773 -788 807 788
<< metal1 >>
rect -813 788 -767 800
rect -813 -788 -807 788
rect -773 -788 -767 788
rect -813 -800 -767 -788
rect -655 788 -609 800
rect -655 -788 -649 788
rect -615 -788 -609 788
rect -655 -800 -609 -788
rect -497 788 -451 800
rect -497 -788 -491 788
rect -457 -788 -451 788
rect -497 -800 -451 -788
rect -339 788 -293 800
rect -339 -788 -333 788
rect -299 -788 -293 788
rect -339 -800 -293 -788
rect -181 788 -135 800
rect -181 -788 -175 788
rect -141 -788 -135 788
rect -181 -800 -135 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 135 788 181 800
rect 135 -788 141 788
rect 175 -788 181 788
rect 135 -800 181 -788
rect 293 788 339 800
rect 293 -788 299 788
rect 333 -788 339 788
rect 293 -800 339 -788
rect 451 788 497 800
rect 451 -788 457 788
rect 491 -788 497 788
rect 451 -800 497 -788
rect 609 788 655 800
rect 609 -788 615 788
rect 649 -788 655 788
rect 609 -800 655 -788
rect 767 788 813 800
rect 767 -788 773 788
rect 807 -788 813 788
rect 767 -800 813 -788
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 0.5 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
