magic
tech sky130A
magscale 1 2
timestamp 1697794495
<< nmos >>
rect -89 -1000 -29 1000
rect 29 -1000 89 1000
<< ndiff >>
rect -147 988 -89 1000
rect -147 -988 -135 988
rect -101 -988 -89 988
rect -147 -1000 -89 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 89 988 147 1000
rect 89 -988 101 988
rect 135 -988 147 988
rect 89 -1000 147 -988
<< ndiffc >>
rect -135 -988 -101 988
rect -17 -988 17 988
rect 101 -988 135 988
<< poly >>
rect -89 1000 -29 1026
rect 29 1000 89 1026
rect -89 -1026 -29 -1000
rect 29 -1026 89 -1000
<< locali >>
rect -135 988 -101 1004
rect -135 -1004 -101 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 101 988 135 1004
rect 101 -1004 135 -988
<< viali >>
rect -135 -988 -101 988
rect -17 -988 17 988
rect 101 -988 135 988
<< metal1 >>
rect -141 988 -95 1000
rect -141 -988 -135 988
rect -101 -988 -95 988
rect -141 -1000 -95 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 95 988 141 1000
rect 95 -988 101 988
rect 135 -988 141 988
rect 95 -1000 141 -988
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 0.3 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
