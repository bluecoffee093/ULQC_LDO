magic
tech sky130A
magscale 1 2
timestamp 1697743316
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
use sky130_fd_pr__nfet_01v8_lvt_Q47UKG  XM1
timestamp 0
transform 1 0 158 0 1 790
box 0 0 1 1
use sky130_fd_pr__pfet_01v8_lvt_AEF6VD  XM2
timestamp 0
transform 1 0 527 0 1 746
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Z
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 A
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 GP
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 GN
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VCCBPIN
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VSSBPIN
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 {}
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 W_N=1
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 L_N=0.35
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 W_P=1
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 L_P=0.35
port 10 nsew
<< end >>
