magic
tech sky130A
magscale 1 2
timestamp 1698954266
<< nwell >>
rect -2571 -299 -2524 -213
rect -918 -299 -872 -212
rect -918 -1340 -873 -1299
rect -2570 -1386 -2455 -1340
rect -987 -1386 -873 -1340
rect 2403 -299 2450 -213
rect 4056 -299 4102 -212
rect 4056 -1340 4101 -1299
rect 2404 -1386 2519 -1340
rect 3987 -1386 4101 -1340
<< pwell >>
rect -228 1435 1760 2076
rect -228 1412 76 1435
rect 1503 1412 1760 1435
rect -228 -2208 1760 1412
rect -2091 -2958 3633 -2208
rect -2091 -2986 -1585 -2958
rect 3117 -2986 3633 -2958
rect -2091 -3304 3633 -2986
rect -2091 -3332 -1585 -3304
rect 3117 -3332 3633 -3304
rect -2091 -4128 3633 -3332
rect -4925 -4571 6548 -4128
rect -4925 -5657 6597 -4571
rect -4925 -11534 6548 -5657
<< psubdiff >>
rect -4974 2086 6597 2120
rect -4974 -4571 -4940 2086
rect -178 1992 1710 2026
rect -178 1379 -144 1992
rect -178 411 -144 1066
rect 1676 1379 1710 1992
rect 1676 411 1710 1066
rect -178 377 1710 411
rect -178 -2258 -144 377
rect 1676 -2258 1710 377
rect -2041 -2292 3583 -2258
rect -2041 -3332 -2007 -2292
rect -2041 -3964 -2007 -3645
rect 3549 -3332 3583 -2292
rect 3549 -3964 3583 -3645
rect -2041 -3998 3583 -3964
rect -4974 -11540 -4940 -5657
rect -4875 -4212 6499 -4178
rect -4875 -4571 -4841 -4212
rect -4875 -11449 -4841 -5657
rect 6465 -4571 6499 -4212
rect 6465 -11449 6499 -5657
rect -4875 -11483 6499 -11449
rect 6563 -4571 6597 2086
rect 6563 -11540 6597 -5657
rect -4974 -11574 6597 -11540
<< psubdiffcont >>
rect -178 1066 -144 1379
rect 1676 1066 1710 1379
rect -2041 -3645 -2007 -3332
rect 3549 -3645 3583 -3332
rect -4974 -5657 -4940 -4571
rect -4875 -5657 -4841 -4571
rect 6465 -5657 6499 -4571
rect 6563 -5657 6597 -4571
<< poly >>
rect 87 1809 1445 1825
rect 87 1806 1103 1809
rect 87 1770 159 1806
rect 193 1770 631 1806
rect 665 1773 1103 1806
rect 1137 1773 1445 1809
rect 665 1770 1445 1773
rect 87 1757 1445 1770
rect 87 1741 147 1757
rect 205 1741 265 1757
rect 323 1741 383 1757
rect 441 1741 501 1757
rect 559 1741 619 1757
rect 677 1741 737 1757
rect 795 1741 855 1757
rect 913 1741 973 1757
rect 1031 1741 1091 1757
rect 1149 1741 1209 1757
rect 1267 1741 1327 1757
rect 1385 1741 1445 1757
rect 87 673 147 689
rect 205 673 265 689
rect 323 673 383 689
rect 441 673 501 689
rect 559 673 619 689
rect 677 673 737 689
rect 795 673 855 689
rect 913 673 973 689
rect 1031 673 1091 689
rect 1149 673 1209 689
rect 1267 673 1327 689
rect 1385 673 1445 689
rect 87 657 1445 673
rect 87 621 159 657
rect 193 621 631 657
rect 665 621 1103 657
rect 1137 621 1445 657
rect 87 605 1445 621
rect -2403 -268 -1039 -202
rect -2403 -1396 -1039 -1330
rect 5 215 105 231
rect 5 85 21 215
rect 89 85 105 215
rect 5 27 105 85
rect 321 189 1211 225
rect 321 105 357 189
rect 1174 105 1211 189
rect 321 69 1211 105
rect 321 27 421 69
rect 479 27 579 69
rect 953 27 1053 69
rect 1111 27 1211 69
rect 1427 215 1527 231
rect 1427 85 1443 215
rect 1511 85 1527 215
rect 1427 27 1527 85
rect 163 -1667 263 -1625
rect 637 -1667 895 -1625
rect 1269 -1667 1369 -1625
rect 163 -1703 1369 -1667
rect 163 -1787 199 -1703
rect 1333 -1787 1369 -1703
rect 163 -1823 1369 -1787
rect 2571 -268 3935 -202
rect 2571 -1396 3935 -1330
rect -1527 -2388 -1327 -2372
rect -1527 -2543 -1511 -2388
rect -1344 -2543 -1327 -2388
rect -1527 -2619 -1327 -2543
rect -1269 -2388 2801 -2372
rect -1269 -2543 -1253 -2388
rect -1085 -2543 -995 -2388
rect -827 -2543 -737 -2388
rect -569 -2543 -479 -2388
rect -311 -2543 -221 -2388
rect -53 -2543 37 -2388
rect 205 -2543 295 -2388
rect 463 -2543 553 -2388
rect 721 -2543 811 -2388
rect 979 -2543 1069 -2388
rect 1237 -2543 1327 -2388
rect 1495 -2543 1585 -2388
rect 1753 -2543 1843 -2388
rect 2011 -2543 2101 -2388
rect 2269 -2543 2359 -2388
rect 2527 -2543 2617 -2388
rect 2785 -2543 2801 -2388
rect -1269 -2598 2801 -2543
rect -1269 -2619 -1069 -2598
rect -1011 -2619 -811 -2598
rect -753 -2619 -553 -2598
rect -495 -2619 -295 -2598
rect -237 -2619 -37 -2598
rect 21 -2619 221 -2598
rect 279 -2619 479 -2598
rect 537 -2619 737 -2598
rect 795 -2619 995 -2598
rect 1053 -2619 1253 -2598
rect 1311 -2619 1511 -2598
rect 1569 -2619 1769 -2598
rect 1827 -2619 2027 -2598
rect 2085 -2619 2285 -2598
rect 2343 -2619 2543 -2598
rect 2601 -2619 2801 -2598
rect 2859 -2388 3059 -2372
rect 2859 -2543 2875 -2388
rect 3043 -2543 3059 -2388
rect 2859 -2619 3059 -2543
rect -1527 -3747 -1327 -3671
rect -1527 -3902 -1511 -3747
rect -1344 -3902 -1327 -3747
rect -1527 -3918 -1327 -3902
rect -1269 -3731 -1069 -3671
rect -1011 -3731 -811 -3671
rect -753 -3731 -553 -3671
rect -495 -3731 -295 -3671
rect -237 -3731 -37 -3671
rect 21 -3731 221 -3671
rect 279 -3731 479 -3671
rect 537 -3731 737 -3671
rect 795 -3731 995 -3671
rect 1053 -3731 1253 -3671
rect 1311 -3731 1511 -3671
rect 1569 -3731 1769 -3671
rect 1827 -3731 2027 -3671
rect 2085 -3731 2285 -3671
rect 2343 -3731 2543 -3671
rect 2601 -3731 2801 -3671
rect -1269 -3747 2801 -3731
rect -1269 -3902 -1253 -3747
rect -1085 -3902 -995 -3747
rect -827 -3902 -737 -3747
rect -569 -3902 -479 -3747
rect -311 -3902 -221 -3747
rect -53 -3902 37 -3747
rect 205 -3902 295 -3747
rect 463 -3902 553 -3747
rect 721 -3902 811 -3747
rect 979 -3902 1069 -3747
rect 1237 -3902 1327 -3747
rect 1495 -3902 1585 -3747
rect 1753 -3902 1843 -3747
rect 2011 -3902 2101 -3747
rect 2269 -3902 2359 -3747
rect 2527 -3902 2617 -3747
rect 2785 -3902 2801 -3747
rect -1269 -3918 2801 -3902
rect 2859 -3747 3059 -3671
rect 2859 -3902 2875 -3747
rect 3043 -3902 3059 -3747
rect 2859 -3918 3059 -3902
<< polycont >>
rect 159 1770 193 1806
rect 631 1770 665 1806
rect 1103 1773 1137 1809
rect 159 621 193 657
rect 631 621 665 657
rect 1103 621 1137 657
rect 21 85 89 215
rect 357 105 1174 189
rect 1443 85 1511 215
rect 199 -1787 1333 -1703
rect -1511 -2543 -1344 -2388
rect -1253 -2543 -1085 -2388
rect -995 -2543 -827 -2388
rect -737 -2543 -569 -2388
rect -479 -2543 -311 -2388
rect -221 -2543 -53 -2388
rect 37 -2543 205 -2388
rect 295 -2543 463 -2388
rect 553 -2543 721 -2388
rect 811 -2543 979 -2388
rect 1069 -2543 1237 -2388
rect 1327 -2543 1495 -2388
rect 1585 -2543 1753 -2388
rect 1843 -2543 2011 -2388
rect 2101 -2543 2269 -2388
rect 2359 -2543 2527 -2388
rect 2617 -2543 2785 -2388
rect 2875 -2543 3043 -2388
rect -1511 -3902 -1344 -3747
rect -1253 -3902 -1085 -3747
rect -995 -3902 -827 -3747
rect -737 -3902 -569 -3747
rect -479 -3902 -311 -3747
rect -221 -3902 -53 -3747
rect 37 -3902 205 -3747
rect 295 -3902 463 -3747
rect 553 -3902 721 -3747
rect 811 -3902 979 -3747
rect 1069 -3902 1237 -3747
rect 1327 -3902 1495 -3747
rect 1585 -3902 1753 -3747
rect 1843 -3902 2011 -3747
rect 2101 -3902 2269 -3747
rect 2359 -3902 2527 -3747
rect 2617 -3902 2785 -3747
rect 2875 -3902 3043 -3747
<< locali >>
rect -4974 2086 6597 2120
rect -4974 -4571 -4940 2086
rect -178 1992 1710 2026
rect -178 1379 -144 1992
rect -178 411 -144 1066
rect 147 1806 205 1825
rect 147 1770 159 1806
rect 193 1770 205 1806
rect 147 657 205 1770
rect 147 621 159 657
rect 193 621 205 657
rect 147 605 205 621
rect 619 1806 677 1825
rect 619 1770 631 1806
rect 665 1770 677 1806
rect 619 657 677 1770
rect 619 621 631 657
rect 665 621 677 657
rect 619 605 677 621
rect 1091 1809 1149 1825
rect 1091 1773 1103 1809
rect 1137 1773 1149 1809
rect 1091 657 1149 1773
rect 1091 621 1103 657
rect 1137 621 1149 657
rect 1091 605 1149 621
rect 1676 1379 1710 1992
rect 1676 411 1710 1066
rect -178 377 1710 411
rect -2678 -1299 -2518 -299
rect -924 -1299 -764 -299
rect -178 -2258 -144 377
rect -53 215 105 231
rect -53 85 21 215
rect 89 85 105 215
rect -53 69 105 85
rect 1427 215 1585 231
rect 1427 85 1443 215
rect 1511 85 1585 215
rect 1427 69 1585 85
rect -53 -1625 5 69
rect 1527 -1625 1585 69
rect 1676 -2258 1710 377
rect 2296 -1299 2456 -299
rect 4050 -1299 4210 -299
rect -2041 -2292 3583 -2258
rect -2041 -3332 -2007 -2292
rect -1573 -2388 -1327 -2372
rect -1573 -2543 -1511 -2388
rect -1344 -2543 -1327 -2388
rect -1573 -2559 -1327 -2543
rect -1269 -2388 2801 -2372
rect -1269 -2543 -1253 -2388
rect -1085 -2394 -995 -2388
rect -827 -2394 -737 -2388
rect -569 -2394 -479 -2388
rect -311 -2394 -221 -2388
rect -53 -2394 37 -2388
rect 205 -2394 295 -2388
rect 463 -2394 553 -2388
rect 721 -2394 811 -2388
rect 979 -2394 1069 -2388
rect 1237 -2394 1327 -2388
rect 1495 -2394 1585 -2388
rect 1753 -2394 1843 -2388
rect 2011 -2394 2101 -2388
rect 2269 -2394 2359 -2388
rect 2527 -2394 2617 -2388
rect -1085 -2543 -995 -2537
rect -827 -2543 -737 -2537
rect -569 -2543 -479 -2537
rect -311 -2543 -221 -2537
rect -53 -2543 37 -2537
rect 205 -2543 295 -2537
rect 463 -2543 553 -2537
rect 721 -2543 811 -2537
rect 979 -2543 1069 -2537
rect 1237 -2543 1327 -2537
rect 1495 -2543 1585 -2537
rect 1753 -2543 1843 -2537
rect 2011 -2543 2101 -2537
rect 2269 -2543 2359 -2537
rect 2527 -2543 2617 -2537
rect 2785 -2543 2801 -2388
rect -1269 -2559 2801 -2543
rect 2859 -2388 3105 -2372
rect 2859 -2543 2875 -2388
rect 3043 -2543 3105 -2388
rect 2859 -2559 3105 -2543
rect -1573 -2641 -1539 -2559
rect 3071 -2641 3105 -2559
rect -1573 -2662 -1539 -2645
rect 3071 -2662 3105 -2645
rect -2041 -3964 -2007 -3645
rect 3549 -3332 3583 -2292
rect -1573 -3731 -1539 -3649
rect 3071 -3731 3105 -3649
rect -1573 -3747 -1327 -3731
rect -1573 -3902 -1511 -3747
rect -1344 -3902 -1327 -3747
rect -1573 -3918 -1327 -3902
rect -1269 -3747 2801 -3731
rect -1269 -3902 -1253 -3747
rect -1085 -3753 -995 -3747
rect -827 -3753 -737 -3747
rect -569 -3753 -479 -3747
rect -311 -3753 -221 -3747
rect -53 -3753 37 -3747
rect 205 -3753 295 -3747
rect 463 -3753 553 -3747
rect 721 -3753 811 -3747
rect 979 -3753 1069 -3747
rect 1237 -3753 1327 -3747
rect 1495 -3753 1585 -3747
rect 1753 -3753 1843 -3747
rect 2011 -3753 2101 -3747
rect 2269 -3753 2359 -3747
rect 2527 -3753 2617 -3747
rect -1085 -3902 -995 -3896
rect -827 -3902 -737 -3896
rect -569 -3902 -479 -3896
rect -311 -3902 -221 -3896
rect -53 -3902 37 -3896
rect 205 -3902 295 -3896
rect 463 -3902 553 -3896
rect 721 -3902 811 -3896
rect 979 -3902 1069 -3896
rect 1237 -3902 1327 -3896
rect 1495 -3902 1585 -3896
rect 1753 -3902 1843 -3896
rect 2011 -3902 2101 -3896
rect 2269 -3902 2359 -3896
rect 2527 -3902 2617 -3896
rect 2785 -3902 2801 -3747
rect -1269 -3918 2801 -3902
rect 2859 -3747 3105 -3731
rect 2859 -3902 2875 -3747
rect 3043 -3902 3105 -3747
rect 2859 -3918 3105 -3902
rect 3549 -3964 3583 -3645
rect -2041 -3998 3583 -3964
rect -4974 -11540 -4940 -5657
rect -4875 -4212 6499 -4178
rect -4875 -4571 -4841 -4212
rect -4875 -11449 -4841 -5657
rect 6465 -4571 6499 -4212
rect 6465 -11449 6499 -5657
rect -4875 -11483 6499 -11449
rect 6563 -4571 6597 2086
rect 6563 -11540 6597 -5657
rect -4974 -11574 6597 -11540
<< viali >>
rect -178 1066 -144 1379
rect 1676 1066 1710 1379
rect 321 189 1211 225
rect 321 105 357 189
rect 357 105 1174 189
rect 1174 105 1211 189
rect 321 69 1211 105
rect 163 -1703 1369 -1667
rect 163 -1787 199 -1703
rect 199 -1787 1333 -1703
rect 1333 -1787 1369 -1703
rect 163 -1823 1369 -1787
rect -1247 -2537 -1085 -2394
rect -1085 -2537 -995 -2394
rect -995 -2537 -827 -2394
rect -827 -2537 -737 -2394
rect -737 -2537 -569 -2394
rect -569 -2537 -479 -2394
rect -479 -2537 -311 -2394
rect -311 -2537 -221 -2394
rect -221 -2537 -53 -2394
rect -53 -2537 37 -2394
rect 37 -2537 205 -2394
rect 205 -2537 295 -2394
rect 295 -2537 463 -2394
rect 463 -2537 553 -2394
rect 553 -2537 721 -2394
rect 721 -2537 811 -2394
rect 811 -2537 979 -2394
rect 979 -2537 1069 -2394
rect 1069 -2537 1237 -2394
rect 1237 -2537 1327 -2394
rect 1327 -2537 1495 -2394
rect 1495 -2537 1585 -2394
rect 1585 -2537 1753 -2394
rect 1753 -2537 1843 -2394
rect 1843 -2537 2011 -2394
rect 2011 -2537 2101 -2394
rect 2101 -2537 2269 -2394
rect 2269 -2537 2359 -2394
rect 2359 -2537 2527 -2394
rect 2527 -2537 2617 -2394
rect 2617 -2537 2779 -2394
rect -2041 -3645 -2007 -3332
rect 3549 -3645 3583 -3332
rect -1247 -3896 -1085 -3753
rect -1085 -3896 -995 -3753
rect -995 -3896 -827 -3753
rect -827 -3896 -737 -3753
rect -737 -3896 -569 -3753
rect -569 -3896 -479 -3753
rect -479 -3896 -311 -3753
rect -311 -3896 -221 -3753
rect -221 -3896 -53 -3753
rect -53 -3896 37 -3753
rect 37 -3896 205 -3753
rect 205 -3896 295 -3753
rect 295 -3896 463 -3753
rect 463 -3896 553 -3753
rect 553 -3896 721 -3753
rect 721 -3896 811 -3753
rect 811 -3896 979 -3753
rect 979 -3896 1069 -3753
rect 1069 -3896 1237 -3753
rect 1237 -3896 1327 -3753
rect 1327 -3896 1495 -3753
rect 1495 -3896 1585 -3753
rect 1585 -3896 1753 -3753
rect 1753 -3896 1843 -3753
rect 1843 -3896 2011 -3753
rect 2011 -3896 2101 -3753
rect 2101 -3896 2269 -3753
rect 2269 -3896 2359 -3753
rect 2359 -3896 2527 -3753
rect 2527 -3896 2617 -3753
rect 2617 -3896 2779 -3753
rect -4974 -5657 -4940 -4571
rect -4875 -5657 -4841 -4571
rect 6465 -5657 6499 -4571
rect 6563 -5657 6597 -4571
<< metal1 >>
rect 29 1391 87 1725
rect -184 1379 87 1391
rect -3203 1369 -2890 1379
rect -3203 1076 -3193 1369
rect -2900 1076 -2890 1369
rect -3203 -3342 -2890 1076
rect -184 1066 -178 1379
rect -144 1366 87 1379
rect -144 1066 29 1366
rect 87 1066 97 1366
rect -184 1054 87 1066
rect 29 715 87 1054
rect 147 1015 205 1825
rect 265 1366 323 1725
rect 383 1715 441 1725
rect 373 1435 383 1715
rect 441 1435 451 1715
rect 255 1066 265 1366
rect 323 1066 333 1366
rect 137 715 147 1015
rect 205 715 215 1015
rect 265 715 323 1066
rect 383 715 441 1435
rect 501 1366 559 1725
rect 491 1066 501 1366
rect 559 1066 569 1366
rect 501 715 559 1066
rect 619 1015 677 1825
rect 737 1366 795 1725
rect 845 1435 855 1715
rect 913 1435 923 1715
rect 727 1066 737 1366
rect 795 1066 805 1366
rect 609 715 619 1015
rect 677 715 687 1015
rect 737 715 795 1066
rect 855 1015 913 1435
rect 973 1366 1031 1725
rect 963 1066 973 1366
rect 1031 1066 1041 1366
rect 973 715 1031 1066
rect 1091 1015 1149 1825
rect 1209 1366 1267 1725
rect 1317 1435 1327 1715
rect 1385 1435 1395 1715
rect 1199 1066 1209 1366
rect 1267 1066 1277 1366
rect 1081 715 1091 1015
rect 1149 715 1159 1015
rect 1209 715 1267 1066
rect 1327 1015 1385 1435
rect 1445 1391 1503 1725
rect 1445 1379 1716 1391
rect 1445 1366 1676 1379
rect 1435 1066 1445 1366
rect 1503 1066 1676 1366
rect 1710 1066 1716 1379
rect 1445 1054 1716 1066
rect 4432 1369 4745 1379
rect 4432 1076 4442 1369
rect 4735 1076 4745 1369
rect 1445 715 1503 1054
rect 147 605 205 715
rect 619 605 677 715
rect 1091 605 1149 715
rect 309 225 1223 231
rect 309 69 321 225
rect 1211 69 1223 225
rect 309 63 1223 69
rect -2688 -268 -2678 -202
rect -2619 -268 -2609 -202
rect -2571 -258 -2455 -212
rect -2678 -649 -2619 -268
rect -2571 -299 -2524 -258
rect -2403 -268 -1039 -202
rect -987 -258 -872 -212
rect -918 -299 -872 -258
rect -833 -268 -823 -202
rect -764 -268 -754 -202
rect -2232 -599 -2222 -299
rect -2164 -599 -2154 -299
rect -1760 -599 -1750 -299
rect -1692 -599 -1682 -299
rect -1288 -599 -1278 -299
rect -1220 -599 -1210 -299
rect -823 -649 -764 -268
rect -53 -527 5 27
rect -2688 -949 -2678 -649
rect -2619 -949 -2609 -649
rect -2468 -949 -2458 -649
rect -2400 -949 -2390 -649
rect -1996 -949 -1986 -649
rect -1928 -949 -1918 -649
rect -1524 -949 -1514 -649
rect -1456 -949 -1446 -649
rect -1052 -949 -1042 -649
rect -984 -949 -974 -649
rect -833 -949 -823 -649
rect -764 -949 -754 -649
rect -2678 -1337 -2619 -949
rect -2586 -1299 -2576 -999
rect -2518 -1299 -2508 -999
rect -2350 -1299 -2340 -999
rect -2282 -1299 -2272 -999
rect -2114 -1299 -2104 -999
rect -2046 -1299 -2036 -999
rect -1878 -1299 -1868 -999
rect -1810 -1299 -1800 -999
rect -1642 -1299 -1632 -999
rect -1574 -1299 -1564 -999
rect -1406 -1299 -1396 -999
rect -1338 -1299 -1328 -999
rect -1170 -1299 -1160 -999
rect -1102 -1299 -1092 -999
rect -934 -1299 -924 -999
rect -866 -1299 -856 -999
rect -2688 -1396 -2678 -1337
rect -2619 -1396 -2609 -1337
rect -2570 -1340 -2524 -1299
rect -2403 -1337 -1039 -1330
rect -2570 -1386 -2455 -1340
rect -2413 -1396 -2403 -1337
rect -1039 -1396 -1029 -1337
rect -918 -1340 -873 -1299
rect -823 -1337 -764 -949
rect -987 -1386 -873 -1340
rect -833 -1396 -823 -1337
rect -764 -1396 -754 -1337
rect -53 -1625 5 -1090
rect 105 -1145 163 1
rect 105 -1625 163 -1599
rect 263 -527 321 27
rect 263 -1625 321 -1090
rect 421 -18 479 8
rect 421 -1625 479 -472
rect 579 -527 637 27
rect 579 -1625 637 -1090
rect 737 -1145 795 1
rect 895 -527 953 27
rect 727 -1599 737 -1145
rect 795 -1599 805 -1145
rect 737 -1625 795 -1599
rect 895 -1625 953 -1090
rect 1053 -18 1111 8
rect 1053 -1625 1111 -472
rect 1211 -527 1269 27
rect 1211 -1625 1269 -1090
rect 1369 -1145 1427 1
rect 1369 -1625 1427 -1599
rect 1527 -527 1585 27
rect 2286 -268 2296 -202
rect 2355 -268 2365 -202
rect 2403 -258 2519 -212
rect 2296 -649 2355 -268
rect 2403 -299 2450 -258
rect 2571 -268 3935 -202
rect 3987 -258 4102 -212
rect 4056 -299 4102 -258
rect 4141 -268 4151 -202
rect 4210 -268 4220 -202
rect 2742 -599 2752 -299
rect 2810 -599 2820 -299
rect 3214 -599 3224 -299
rect 3282 -599 3292 -299
rect 3686 -599 3696 -299
rect 3754 -599 3764 -299
rect 4151 -649 4210 -268
rect 2286 -949 2296 -649
rect 2355 -949 2365 -649
rect 2506 -949 2516 -649
rect 2574 -949 2584 -649
rect 2978 -949 2988 -649
rect 3046 -949 3056 -649
rect 3450 -949 3460 -649
rect 3518 -949 3528 -649
rect 3922 -949 3932 -649
rect 3990 -949 4000 -649
rect 4141 -949 4151 -649
rect 4210 -949 4220 -649
rect 1527 -1625 1585 -1090
rect 2296 -1337 2355 -949
rect 2388 -1299 2398 -999
rect 2456 -1299 2466 -999
rect 2624 -1299 2634 -999
rect 2692 -1299 2702 -999
rect 2860 -1299 2870 -999
rect 2928 -1299 2938 -999
rect 3096 -1299 3106 -999
rect 3164 -1299 3174 -999
rect 3332 -1299 3342 -999
rect 3400 -1299 3410 -999
rect 3568 -1299 3578 -999
rect 3636 -1299 3646 -999
rect 3804 -1299 3814 -999
rect 3872 -1299 3882 -999
rect 4040 -1299 4050 -999
rect 4108 -1299 4118 -999
rect 2286 -1396 2296 -1337
rect 2355 -1396 2365 -1337
rect 2404 -1340 2450 -1299
rect 2571 -1337 3935 -1330
rect 2404 -1386 2519 -1340
rect 2561 -1396 2571 -1337
rect 3935 -1396 3945 -1337
rect 4056 -1340 4101 -1299
rect 4151 -1337 4210 -949
rect 3987 -1386 4101 -1340
rect 4141 -1396 4151 -1337
rect 4210 -1396 4220 -1337
rect 151 -1667 1381 -1661
rect 151 -1823 163 -1667
rect 1369 -1823 1381 -1667
rect 151 -1829 1381 -1823
rect -1942 -2382 -1697 -2372
rect -1942 -2597 -1932 -2382
rect -1707 -2597 -1697 -2382
rect -1942 -2996 -1697 -2597
rect -1269 -2607 -1259 -2382
rect 2791 -2607 2801 -2382
rect 3239 -2388 3484 -2372
rect 3239 -2603 3249 -2388
rect 3474 -2603 3484 -2388
rect -1337 -2948 -1327 -2655
rect -1269 -2948 -1259 -2655
rect -305 -2948 -295 -2655
rect -237 -2948 -227 -2655
rect 727 -2948 737 -2655
rect 795 -2948 805 -2655
rect 1759 -2948 1769 -2655
rect 1827 -2948 1837 -2655
rect 2791 -2948 2801 -2655
rect 2859 -2948 2869 -2655
rect 3239 -2996 3484 -2603
rect -1942 -3294 -1932 -2996
rect -1707 -3294 -1697 -2996
rect -821 -3294 -811 -2996
rect -753 -3294 -743 -2996
rect 211 -3294 221 -2996
rect 279 -3294 289 -2996
rect 1243 -3294 1253 -2996
rect 1311 -3294 1321 -2996
rect 2275 -3294 2285 -2996
rect 2343 -3294 2353 -2996
rect 3239 -3294 3249 -2996
rect 3474 -3294 3484 -2996
rect -3203 -3635 -3193 -3342
rect -2900 -3635 -2890 -3342
rect -3203 -3645 -2890 -3635
rect -2091 -3332 -2001 -3320
rect -2091 -3657 -2001 -3645
rect -1942 -3683 -1697 -3294
rect -1595 -3635 -1585 -3342
rect -1527 -3635 -1517 -3342
rect -1079 -3635 -1069 -3342
rect -1011 -3635 -1001 -3342
rect -563 -3635 -553 -3342
rect -495 -3635 -485 -3342
rect -47 -3635 -37 -3342
rect 21 -3635 31 -3342
rect 469 -3635 479 -3342
rect 537 -3635 547 -3342
rect 985 -3635 995 -3342
rect 1053 -3635 1063 -3342
rect 1501 -3635 1511 -3342
rect 1569 -3635 1579 -3342
rect 2017 -3635 2027 -3342
rect 2085 -3635 2095 -3342
rect 2533 -3635 2543 -3342
rect 2601 -3635 2611 -3342
rect 3049 -3635 3059 -3342
rect 3117 -3635 3127 -3342
rect -1942 -3908 -1932 -3683
rect -1707 -3908 -1697 -3683
rect -1942 -3918 -1697 -3908
rect -1269 -3683 2801 -3673
rect -1269 -3908 -1259 -3683
rect 2791 -3908 2801 -3683
rect -1269 -3918 2801 -3908
rect 3239 -3693 3484 -3294
rect 3543 -3332 3633 -3320
rect 4432 -3342 4745 1076
rect 4432 -3635 4442 -3342
rect 4735 -3635 4745 -3342
rect 4432 -3645 4745 -3635
rect 3543 -3657 3633 -3645
rect 3239 -3908 3249 -3693
rect 3474 -3908 3484 -3693
rect 3239 -3918 3484 -3908
rect -4801 -4435 -4791 -4262
rect -4584 -4435 -4574 -4262
rect 6198 -4435 6208 -4262
rect 6415 -4435 6425 -4262
rect -4980 -4571 -4934 -4559
rect -4881 -4571 -4835 -4559
rect -4984 -5657 -4974 -4571
rect -4841 -5657 -4831 -4571
rect -4980 -5669 -4934 -5657
rect -4881 -5669 -4835 -5657
rect -4791 -5853 -4584 -4435
rect 6208 -4571 6415 -4435
rect 6459 -4571 6505 -4559
rect 6557 -4571 6603 -4559
rect -4375 -4745 -4365 -4571
rect -4159 -4745 -4149 -4571
rect -3933 -4735 -3923 -4679
rect -3857 -4735 -3847 -4679
rect -3741 -4735 -3731 -4679
rect -3665 -4735 -3655 -4679
rect -3549 -4735 -3539 -4679
rect -3473 -4735 -3463 -4679
rect -3357 -4735 -3347 -4679
rect -3281 -4735 -3271 -4679
rect -3165 -4735 -3155 -4679
rect -3089 -4735 -3079 -4679
rect -2973 -4735 -2963 -4679
rect -2897 -4735 -2887 -4679
rect -2781 -4735 -2771 -4679
rect -2705 -4735 -2695 -4679
rect -2589 -4735 -2579 -4679
rect -2513 -4735 -2503 -4679
rect -2397 -4735 -2387 -4679
rect -2321 -4735 -2311 -4679
rect -2205 -4735 -2195 -4679
rect -2129 -4735 -2119 -4679
rect -2013 -4735 -2003 -4679
rect -1937 -4735 -1927 -4679
rect -1821 -4735 -1811 -4679
rect -1745 -4735 -1735 -4679
rect -1629 -4735 -1619 -4679
rect -1553 -4735 -1543 -4679
rect -1437 -4735 -1427 -4679
rect -1361 -4735 -1351 -4679
rect -1245 -4735 -1235 -4679
rect -1169 -4735 -1159 -4679
rect -1053 -4735 -1043 -4679
rect -977 -4735 -967 -4679
rect -861 -4735 -851 -4679
rect -785 -4735 -775 -4679
rect -669 -4735 -659 -4679
rect -593 -4735 -583 -4679
rect -477 -4735 -467 -4679
rect -401 -4735 -391 -4679
rect -285 -4735 -275 -4679
rect -209 -4735 -199 -4679
rect -93 -4735 -83 -4679
rect -17 -4735 -7 -4679
rect 99 -4735 109 -4679
rect 175 -4735 185 -4679
rect 291 -4735 301 -4679
rect 367 -4735 377 -4679
rect 483 -4735 493 -4679
rect 559 -4735 569 -4679
rect 675 -4735 685 -4679
rect 751 -4735 761 -4679
rect 867 -4735 877 -4679
rect 943 -4735 953 -4679
rect 1059 -4735 1069 -4679
rect 1135 -4735 1145 -4679
rect 1251 -4735 1261 -4679
rect 1327 -4735 1337 -4679
rect 1443 -4735 1453 -4679
rect 1519 -4735 1529 -4679
rect 1635 -4735 1645 -4679
rect 1711 -4735 1721 -4679
rect 1827 -4735 1837 -4679
rect 1903 -4735 1913 -4679
rect 2019 -4735 2029 -4679
rect 2095 -4735 2105 -4679
rect 2211 -4735 2221 -4679
rect 2287 -4735 2297 -4679
rect 2403 -4735 2413 -4679
rect 2479 -4735 2489 -4679
rect 2595 -4735 2605 -4679
rect 2671 -4735 2681 -4679
rect 2787 -4735 2797 -4679
rect 2863 -4735 2873 -4679
rect 2979 -4735 2989 -4679
rect 3055 -4735 3065 -4679
rect 3171 -4735 3181 -4679
rect 3247 -4735 3257 -4679
rect 3363 -4735 3373 -4679
rect 3439 -4735 3449 -4679
rect 3555 -4735 3565 -4679
rect 3631 -4735 3641 -4679
rect 3747 -4735 3757 -4679
rect 3823 -4735 3833 -4679
rect 3939 -4735 3949 -4679
rect 4015 -4735 4025 -4679
rect 4131 -4735 4141 -4679
rect 4207 -4735 4217 -4679
rect 4323 -4735 4333 -4679
rect 4399 -4735 4409 -4679
rect 4515 -4735 4525 -4679
rect 4591 -4735 4601 -4679
rect 4707 -4735 4717 -4679
rect 4783 -4735 4793 -4679
rect 4899 -4735 4909 -4679
rect 4975 -4735 4985 -4679
rect 5091 -4735 5101 -4679
rect 5167 -4735 5177 -4679
rect 5283 -4735 5293 -4679
rect 5359 -4735 5369 -4679
rect 5475 -4735 5485 -4679
rect 5551 -4735 5561 -4679
rect 5681 -4745 5691 -4571
rect 5897 -4745 5907 -4571
rect -4365 -4956 -4159 -4745
rect -4063 -4956 -4011 -4950
rect -4375 -5657 -4365 -4956
rect -4159 -5657 -4149 -4956
rect -4800 -6564 -4790 -5853
rect -4584 -6564 -4574 -5853
rect -4791 -8071 -4584 -6564
rect -4365 -6789 -4159 -5657
rect -4063 -5664 -4011 -5657
rect -3871 -4956 -3819 -4950
rect -3871 -5664 -3819 -5657
rect -3679 -4956 -3627 -4950
rect -3679 -5664 -3627 -5657
rect -3487 -4956 -3435 -4950
rect -3487 -5664 -3435 -5657
rect -3295 -4956 -3243 -4950
rect -3295 -5664 -3243 -5657
rect -3103 -4956 -3051 -4950
rect -3103 -5664 -3051 -5657
rect -2911 -4956 -2859 -4950
rect -2911 -5664 -2859 -5657
rect -2719 -4956 -2667 -4950
rect -2719 -5664 -2667 -5657
rect -2527 -4956 -2475 -4950
rect -2527 -5664 -2475 -5657
rect -2335 -4956 -2283 -4950
rect -2335 -5664 -2283 -5657
rect -2143 -4956 -2091 -4950
rect -2143 -5664 -2091 -5657
rect -1951 -4956 -1899 -4950
rect -1951 -5664 -1899 -5657
rect -1759 -4956 -1707 -4950
rect -1759 -5664 -1707 -5657
rect -1567 -4956 -1515 -4950
rect -1567 -5664 -1515 -5657
rect -1375 -4956 -1323 -4950
rect -1375 -5664 -1323 -5657
rect -1183 -4956 -1131 -4950
rect -1183 -5664 -1131 -5657
rect -991 -4956 -939 -4950
rect -991 -5664 -939 -5657
rect -799 -4956 -747 -4950
rect -799 -5664 -747 -5657
rect -607 -4956 -555 -4950
rect -607 -5664 -555 -5657
rect -415 -4956 -363 -4950
rect -415 -5664 -363 -5657
rect -223 -4956 -171 -4950
rect -223 -5664 -171 -5657
rect -31 -4956 21 -4950
rect -31 -5664 21 -5657
rect 161 -4956 213 -4950
rect 161 -5664 213 -5657
rect 353 -4956 405 -4950
rect 353 -5664 405 -5657
rect 545 -4956 597 -4950
rect 545 -5664 597 -5657
rect 737 -4956 789 -4950
rect 737 -5664 789 -5657
rect 929 -4956 981 -4950
rect 929 -5664 981 -5657
rect 1121 -4956 1173 -4950
rect 1121 -5664 1173 -5657
rect 1313 -4956 1365 -4950
rect 1313 -5664 1365 -5657
rect 1505 -4956 1557 -4950
rect 1505 -5664 1557 -5657
rect 1697 -4956 1749 -4950
rect 1697 -5664 1749 -5657
rect 1889 -4956 1941 -4950
rect 1889 -5664 1941 -5657
rect 2081 -4956 2133 -4950
rect 2081 -5664 2133 -5657
rect 2273 -4956 2325 -4950
rect 2273 -5664 2325 -5657
rect 2465 -4956 2517 -4950
rect 2465 -5664 2517 -5657
rect 2657 -4956 2709 -4950
rect 2657 -5664 2709 -5657
rect 2849 -4956 2901 -4950
rect 2849 -5664 2901 -5657
rect 3041 -4956 3093 -4950
rect 3041 -5664 3093 -5657
rect 3233 -4956 3285 -4950
rect 3233 -5664 3285 -5657
rect 3425 -4956 3477 -4950
rect 3425 -5664 3477 -5657
rect 3617 -4956 3669 -4950
rect 3617 -5664 3669 -5657
rect 3809 -4956 3861 -4950
rect 3809 -5664 3861 -5657
rect 4001 -4956 4053 -4950
rect 4001 -5664 4053 -5657
rect 4193 -4956 4245 -4950
rect 4193 -5664 4245 -5657
rect 4385 -4956 4437 -4950
rect 4385 -5664 4437 -5657
rect 4577 -4956 4629 -4950
rect 4577 -5664 4629 -5657
rect 4769 -4956 4821 -4950
rect 4769 -5664 4821 -5657
rect 4961 -4956 5013 -4950
rect 4961 -5664 5013 -5657
rect 5153 -4956 5205 -4950
rect 5153 -5664 5205 -5657
rect 5345 -4956 5397 -4950
rect 5691 -4956 5897 -4745
rect 5527 -5657 5537 -4956
rect 5589 -5657 5599 -4956
rect 5681 -5657 5691 -4956
rect 5897 -5657 5907 -4956
rect 5345 -5664 5397 -5657
rect -3971 -5853 -3905 -5843
rect -3971 -6574 -3905 -6564
rect -3779 -5853 -3713 -5843
rect -3779 -6574 -3713 -6564
rect -3587 -5853 -3521 -5843
rect -3587 -6574 -3521 -6564
rect -3395 -5853 -3329 -5843
rect -3395 -6574 -3329 -6564
rect -3203 -5853 -3137 -5843
rect -3203 -6574 -3137 -6564
rect -3011 -5853 -2945 -5843
rect -3011 -6574 -2945 -6564
rect -2819 -5853 -2753 -5843
rect -2819 -6574 -2753 -6564
rect -2627 -5853 -2561 -5843
rect -2627 -6574 -2561 -6564
rect -2435 -5853 -2369 -5843
rect -2435 -6574 -2369 -6564
rect -2243 -5853 -2177 -5843
rect -2243 -6574 -2177 -6564
rect -2051 -5853 -1985 -5843
rect -2051 -6574 -1985 -6564
rect -1859 -5853 -1793 -5843
rect -1859 -6574 -1793 -6564
rect -1667 -5853 -1601 -5843
rect -1667 -6574 -1601 -6564
rect -1475 -5853 -1409 -5843
rect -1475 -6574 -1409 -6564
rect -1283 -5853 -1217 -5843
rect -1283 -6574 -1217 -6564
rect -1091 -5853 -1025 -5843
rect -1091 -6574 -1025 -6564
rect -899 -5853 -833 -5843
rect -899 -6574 -833 -6564
rect -707 -5853 -641 -5843
rect -707 -6574 -641 -6564
rect -515 -5853 -449 -5843
rect -515 -6574 -449 -6564
rect -323 -5853 -257 -5843
rect -323 -6574 -257 -6564
rect -131 -5853 -65 -5843
rect -131 -6574 -65 -6564
rect 61 -5853 127 -5843
rect 61 -6574 127 -6564
rect 253 -5853 319 -5843
rect 253 -6574 319 -6564
rect 445 -5853 511 -5843
rect 445 -6574 511 -6564
rect 637 -5853 703 -5843
rect 637 -6574 703 -6564
rect 829 -5853 895 -5843
rect 829 -6574 895 -6564
rect 1021 -5853 1087 -5843
rect 1021 -6574 1087 -6564
rect 1213 -5853 1279 -5843
rect 1213 -6574 1279 -6564
rect 1405 -5853 1471 -5843
rect 1405 -6574 1471 -6564
rect 1597 -5853 1663 -5843
rect 1597 -6574 1663 -6564
rect 1789 -5853 1855 -5843
rect 1789 -6574 1855 -6564
rect 1981 -5853 2047 -5843
rect 1981 -6574 2047 -6564
rect 2173 -5853 2239 -5843
rect 2173 -6574 2239 -6564
rect 2365 -5853 2431 -5843
rect 2365 -6574 2431 -6564
rect 2557 -5853 2623 -5843
rect 2557 -6574 2623 -6564
rect 2749 -5853 2815 -5843
rect 2749 -6574 2815 -6564
rect 2941 -5853 3007 -5843
rect 2941 -6574 3007 -6564
rect 3133 -5853 3199 -5843
rect 3133 -6574 3199 -6564
rect 3325 -5853 3391 -5843
rect 3325 -6574 3391 -6564
rect 3517 -5853 3583 -5843
rect 3517 -6574 3583 -6564
rect 3709 -5853 3775 -5843
rect 3709 -6574 3775 -6564
rect 3901 -5853 3967 -5843
rect 3901 -6574 3967 -6564
rect 4093 -5853 4159 -5843
rect 4093 -6574 4159 -6564
rect 4285 -5853 4351 -5843
rect 4285 -6574 4351 -6564
rect 4477 -5853 4543 -5843
rect 4477 -6574 4543 -6564
rect 4669 -5853 4735 -5843
rect 4669 -6574 4735 -6564
rect 4861 -5853 4927 -5843
rect 4861 -6574 4927 -6564
rect 5053 -5853 5119 -5843
rect 5053 -6574 5119 -6564
rect 5245 -5853 5311 -5843
rect 5245 -6574 5311 -6564
rect 5437 -5853 5503 -5843
rect 5437 -6574 5503 -6564
rect 5691 -6789 5897 -5657
rect 6208 -5853 6414 -4571
rect 6455 -5657 6465 -4571
rect 6598 -5657 6608 -4571
rect 6459 -5669 6505 -5657
rect 6557 -5669 6603 -5657
rect 6198 -6564 6208 -5853
rect 6414 -6564 6424 -5853
rect -4375 -6963 -4365 -6789
rect -4159 -6963 -4149 -6789
rect -4029 -6855 -4019 -6799
rect -3953 -6855 -3943 -6799
rect -3837 -6855 -3827 -6799
rect -3761 -6855 -3751 -6799
rect -3645 -6855 -3635 -6799
rect -3569 -6855 -3559 -6799
rect -3453 -6855 -3443 -6799
rect -3377 -6855 -3367 -6799
rect -3261 -6855 -3251 -6799
rect -3185 -6855 -3175 -6799
rect -3069 -6855 -3059 -6799
rect -2993 -6855 -2983 -6799
rect -2877 -6855 -2867 -6799
rect -2801 -6855 -2791 -6799
rect -2685 -6855 -2675 -6799
rect -2609 -6855 -2599 -6799
rect -2493 -6855 -2483 -6799
rect -2417 -6855 -2407 -6799
rect -2301 -6855 -2291 -6799
rect -2225 -6855 -2215 -6799
rect -2109 -6855 -2099 -6799
rect -2033 -6855 -2023 -6799
rect -1917 -6855 -1907 -6799
rect -1841 -6855 -1831 -6799
rect -1725 -6855 -1715 -6799
rect -1649 -6855 -1639 -6799
rect -1533 -6855 -1523 -6799
rect -1457 -6855 -1447 -6799
rect -1341 -6855 -1331 -6799
rect -1265 -6855 -1255 -6799
rect -1149 -6855 -1139 -6799
rect -1073 -6855 -1063 -6799
rect -957 -6855 -947 -6799
rect -881 -6855 -871 -6799
rect -765 -6855 -755 -6799
rect -689 -6855 -679 -6799
rect -573 -6855 -563 -6799
rect -497 -6855 -487 -6799
rect -381 -6855 -371 -6799
rect -305 -6855 -295 -6799
rect -189 -6855 -179 -6799
rect -113 -6855 -103 -6799
rect 3 -6855 13 -6799
rect 79 -6855 89 -6799
rect 195 -6855 205 -6799
rect 271 -6855 281 -6799
rect 387 -6855 397 -6799
rect 463 -6855 473 -6799
rect 579 -6855 589 -6799
rect 655 -6855 665 -6799
rect 771 -6855 781 -6799
rect 847 -6855 857 -6799
rect 963 -6855 973 -6799
rect 1039 -6855 1049 -6799
rect 1155 -6855 1165 -6799
rect 1231 -6855 1241 -6799
rect 1347 -6855 1357 -6799
rect 1423 -6855 1433 -6799
rect 1539 -6855 1549 -6799
rect 1615 -6855 1625 -6799
rect 1731 -6855 1741 -6799
rect 1807 -6855 1817 -6799
rect 1923 -6855 1933 -6799
rect 1999 -6855 2009 -6799
rect 2115 -6855 2125 -6799
rect 2191 -6855 2201 -6799
rect 2307 -6855 2317 -6799
rect 2383 -6855 2393 -6799
rect 2499 -6855 2509 -6799
rect 2575 -6855 2585 -6799
rect 2691 -6855 2701 -6799
rect 2767 -6855 2777 -6799
rect 2883 -6855 2893 -6799
rect 2959 -6855 2969 -6799
rect 3075 -6855 3085 -6799
rect 3151 -6855 3161 -6799
rect 3267 -6855 3277 -6799
rect 3343 -6855 3353 -6799
rect 3459 -6855 3469 -6799
rect 3535 -6855 3545 -6799
rect 3651 -6855 3661 -6799
rect 3727 -6855 3737 -6799
rect 3843 -6855 3853 -6799
rect 3919 -6855 3929 -6799
rect 4035 -6855 4045 -6799
rect 4111 -6855 4121 -6799
rect 4227 -6855 4237 -6799
rect 4303 -6855 4313 -6799
rect 4419 -6855 4429 -6799
rect 4495 -6855 4505 -6799
rect 4611 -6855 4621 -6799
rect 4687 -6855 4697 -6799
rect 4803 -6855 4813 -6799
rect 4879 -6855 4889 -6799
rect 4995 -6855 5005 -6799
rect 5071 -6855 5081 -6799
rect 5187 -6855 5197 -6799
rect 5263 -6855 5273 -6799
rect 5379 -6855 5389 -6799
rect 5455 -6855 5465 -6799
rect -4029 -6953 -4019 -6897
rect -3953 -6953 -3943 -6897
rect -3837 -6953 -3827 -6897
rect -3761 -6953 -3751 -6897
rect -3645 -6953 -3635 -6897
rect -3569 -6953 -3559 -6897
rect -3453 -6953 -3443 -6897
rect -3377 -6953 -3367 -6897
rect -3261 -6953 -3251 -6897
rect -3185 -6953 -3175 -6897
rect -3069 -6953 -3059 -6897
rect -2993 -6953 -2983 -6897
rect -2877 -6953 -2867 -6897
rect -2801 -6953 -2791 -6897
rect -2685 -6953 -2675 -6897
rect -2609 -6953 -2599 -6897
rect -2493 -6953 -2483 -6897
rect -2417 -6953 -2407 -6897
rect -2301 -6953 -2291 -6897
rect -2225 -6953 -2215 -6897
rect -2109 -6953 -2099 -6897
rect -2033 -6953 -2023 -6897
rect -1917 -6953 -1907 -6897
rect -1841 -6953 -1831 -6897
rect -1725 -6953 -1715 -6897
rect -1649 -6953 -1639 -6897
rect -1533 -6953 -1523 -6897
rect -1457 -6953 -1447 -6897
rect -1341 -6953 -1331 -6897
rect -1265 -6953 -1255 -6897
rect -1149 -6953 -1139 -6897
rect -1073 -6953 -1063 -6897
rect -957 -6953 -947 -6897
rect -881 -6953 -871 -6897
rect -765 -6953 -755 -6897
rect -689 -6953 -679 -6897
rect -573 -6953 -563 -6897
rect -497 -6953 -487 -6897
rect -381 -6953 -371 -6897
rect -305 -6953 -295 -6897
rect -189 -6953 -179 -6897
rect -113 -6953 -103 -6897
rect 3 -6953 13 -6897
rect 79 -6953 89 -6897
rect 195 -6953 205 -6897
rect 271 -6953 281 -6897
rect 387 -6953 397 -6897
rect 463 -6953 473 -6897
rect 579 -6953 589 -6897
rect 655 -6953 665 -6897
rect 771 -6953 781 -6897
rect 847 -6953 857 -6897
rect 963 -6953 973 -6897
rect 1039 -6953 1049 -6897
rect 1155 -6953 1165 -6897
rect 1231 -6953 1241 -6897
rect 1347 -6953 1357 -6897
rect 1423 -6953 1433 -6897
rect 1539 -6953 1549 -6897
rect 1615 -6953 1625 -6897
rect 1731 -6953 1741 -6897
rect 1807 -6953 1817 -6897
rect 1923 -6953 1933 -6897
rect 1999 -6953 2009 -6897
rect 2115 -6953 2125 -6897
rect 2191 -6953 2201 -6897
rect 2307 -6953 2317 -6897
rect 2383 -6953 2393 -6897
rect 2499 -6953 2509 -6897
rect 2575 -6953 2585 -6897
rect 2691 -6953 2701 -6897
rect 2767 -6953 2777 -6897
rect 2883 -6953 2893 -6897
rect 2959 -6953 2969 -6897
rect 3075 -6953 3085 -6897
rect 3151 -6953 3161 -6897
rect 3267 -6953 3277 -6897
rect 3343 -6953 3353 -6897
rect 3459 -6953 3469 -6897
rect 3535 -6953 3545 -6897
rect 3651 -6953 3661 -6897
rect 3727 -6953 3737 -6897
rect 3843 -6953 3853 -6897
rect 3919 -6953 3929 -6897
rect 4035 -6953 4045 -6897
rect 4111 -6953 4121 -6897
rect 4227 -6953 4237 -6897
rect 4303 -6953 4313 -6897
rect 4419 -6953 4429 -6897
rect 4495 -6953 4505 -6897
rect 4611 -6953 4621 -6897
rect 4687 -6953 4697 -6897
rect 4803 -6953 4813 -6897
rect 4879 -6953 4889 -6897
rect 4995 -6953 5005 -6897
rect 5071 -6953 5081 -6897
rect 5187 -6953 5197 -6897
rect 5263 -6953 5273 -6897
rect 5379 -6953 5389 -6897
rect 5455 -6953 5465 -6897
rect 5681 -6963 5691 -6789
rect 5897 -6963 5907 -6789
rect -4365 -7174 -4159 -6963
rect -4063 -7174 -4011 -7164
rect -4375 -7875 -4365 -7174
rect -4159 -7875 -4149 -7174
rect -4800 -8782 -4790 -8071
rect -4584 -8782 -4574 -8071
rect -4791 -10289 -4584 -8782
rect -4365 -9007 -4159 -7875
rect -4063 -7885 -4011 -7875
rect -3871 -7174 -3819 -7164
rect -3871 -7885 -3819 -7875
rect -3679 -7174 -3627 -7164
rect -3679 -7885 -3627 -7875
rect -3487 -7174 -3435 -7164
rect -3487 -7885 -3435 -7875
rect -3295 -7174 -3243 -7164
rect -3295 -7885 -3243 -7875
rect -3103 -7174 -3051 -7164
rect -3103 -7885 -3051 -7875
rect -2911 -7174 -2859 -7164
rect -2911 -7885 -2859 -7875
rect -2719 -7174 -2667 -7164
rect -2719 -7885 -2667 -7875
rect -2527 -7174 -2475 -7164
rect -2527 -7885 -2475 -7875
rect -2335 -7174 -2283 -7164
rect -2335 -7885 -2283 -7875
rect -2143 -7174 -2091 -7164
rect -2143 -7885 -2091 -7875
rect -1951 -7174 -1899 -7164
rect -1951 -7885 -1899 -7875
rect -1759 -7174 -1707 -7164
rect -1759 -7885 -1707 -7875
rect -1567 -7174 -1515 -7164
rect -1567 -7885 -1515 -7875
rect -1375 -7174 -1323 -7164
rect -1375 -7885 -1323 -7875
rect -1183 -7174 -1131 -7164
rect -1183 -7885 -1131 -7875
rect -991 -7174 -939 -7164
rect -991 -7885 -939 -7875
rect -799 -7174 -747 -7164
rect -799 -7885 -747 -7875
rect -607 -7174 -555 -7164
rect -607 -7885 -555 -7875
rect -415 -7174 -363 -7164
rect -415 -7885 -363 -7875
rect -223 -7174 -171 -7164
rect -223 -7885 -171 -7875
rect -31 -7174 21 -7164
rect -31 -7885 21 -7875
rect 161 -7174 213 -7164
rect 161 -7885 213 -7875
rect 353 -7174 405 -7164
rect 353 -7885 405 -7875
rect 545 -7174 597 -7164
rect 545 -7885 597 -7875
rect 737 -7174 789 -7164
rect 737 -7885 789 -7875
rect 929 -7174 981 -7164
rect 929 -7885 981 -7875
rect 1121 -7174 1173 -7164
rect 1121 -7885 1173 -7875
rect 1313 -7174 1365 -7164
rect 1313 -7885 1365 -7875
rect 1505 -7174 1557 -7164
rect 1505 -7885 1557 -7875
rect 1697 -7174 1749 -7164
rect 1697 -7885 1749 -7875
rect 1889 -7174 1941 -7164
rect 1889 -7885 1941 -7875
rect 2081 -7174 2133 -7164
rect 2081 -7885 2133 -7875
rect 2273 -7174 2325 -7164
rect 2273 -7885 2325 -7875
rect 2465 -7174 2517 -7164
rect 2465 -7885 2517 -7875
rect 2657 -7174 2709 -7164
rect 2657 -7885 2709 -7875
rect 2849 -7174 2901 -7164
rect 2849 -7885 2901 -7875
rect 3041 -7174 3093 -7164
rect 3041 -7885 3093 -7875
rect 3233 -7174 3285 -7164
rect 3233 -7885 3285 -7875
rect 3425 -7174 3477 -7164
rect 3425 -7885 3477 -7875
rect 3617 -7174 3669 -7164
rect 3617 -7885 3669 -7875
rect 3809 -7174 3861 -7164
rect 3809 -7885 3861 -7875
rect 4001 -7174 4053 -7164
rect 4001 -7885 4053 -7875
rect 4193 -7174 4245 -7164
rect 4193 -7885 4245 -7875
rect 4385 -7174 4437 -7164
rect 4385 -7885 4437 -7875
rect 4577 -7174 4629 -7164
rect 4577 -7885 4629 -7875
rect 4769 -7174 4821 -7164
rect 4769 -7885 4821 -7875
rect 4961 -7174 5013 -7164
rect 4961 -7885 5013 -7875
rect 5153 -7174 5205 -7164
rect 5153 -7885 5205 -7875
rect 5345 -7174 5397 -7164
rect 5691 -7174 5897 -6963
rect 5527 -7875 5537 -7174
rect 5589 -7875 5599 -7174
rect 5681 -7875 5691 -7174
rect 5897 -7875 5907 -7174
rect 5345 -7885 5397 -7875
rect -3971 -8071 -3905 -8061
rect -3971 -8792 -3905 -8782
rect -3779 -8071 -3713 -8061
rect -3779 -8792 -3713 -8782
rect -3587 -8071 -3521 -8061
rect -3587 -8792 -3521 -8782
rect -3395 -8071 -3329 -8061
rect -3395 -8792 -3329 -8782
rect -3203 -8071 -3137 -8061
rect -3203 -8792 -3137 -8782
rect -3011 -8071 -2945 -8061
rect -3011 -8792 -2945 -8782
rect -2819 -8071 -2753 -8061
rect -2819 -8792 -2753 -8782
rect -2627 -8071 -2561 -8061
rect -2627 -8792 -2561 -8782
rect -2435 -8071 -2369 -8061
rect -2435 -8792 -2369 -8782
rect -2243 -8071 -2177 -8061
rect -2243 -8792 -2177 -8782
rect -2051 -8071 -1985 -8061
rect -2051 -8792 -1985 -8782
rect -1859 -8071 -1793 -8061
rect -1859 -8792 -1793 -8782
rect -1667 -8071 -1601 -8061
rect -1667 -8792 -1601 -8782
rect -1475 -8071 -1409 -8061
rect -1475 -8792 -1409 -8782
rect -1283 -8071 -1217 -8061
rect -1283 -8792 -1217 -8782
rect -1091 -8071 -1025 -8061
rect -1091 -8792 -1025 -8782
rect -899 -8071 -833 -8061
rect -899 -8792 -833 -8782
rect -707 -8071 -641 -8061
rect -707 -8792 -641 -8782
rect -515 -8071 -449 -8061
rect -515 -8792 -449 -8782
rect -323 -8071 -257 -8061
rect -323 -8792 -257 -8782
rect -131 -8071 -65 -8061
rect -131 -8792 -65 -8782
rect 61 -8071 127 -8061
rect 61 -8792 127 -8782
rect 253 -8071 319 -8061
rect 253 -8792 319 -8782
rect 445 -8071 511 -8061
rect 445 -8792 511 -8782
rect 637 -8071 703 -8061
rect 637 -8792 703 -8782
rect 829 -8071 895 -8061
rect 829 -8792 895 -8782
rect 1021 -8071 1087 -8061
rect 1021 -8792 1087 -8782
rect 1213 -8071 1279 -8061
rect 1213 -8792 1279 -8782
rect 1405 -8071 1471 -8061
rect 1405 -8792 1471 -8782
rect 1597 -8071 1663 -8061
rect 1597 -8792 1663 -8782
rect 1789 -8071 1855 -8061
rect 1789 -8792 1855 -8782
rect 1981 -8071 2047 -8061
rect 1981 -8792 2047 -8782
rect 2173 -8071 2239 -8061
rect 2173 -8792 2239 -8782
rect 2365 -8071 2431 -8061
rect 2365 -8792 2431 -8782
rect 2557 -8071 2623 -8061
rect 2557 -8792 2623 -8782
rect 2749 -8071 2815 -8061
rect 2749 -8792 2815 -8782
rect 2941 -8071 3007 -8061
rect 2941 -8792 3007 -8782
rect 3133 -8071 3199 -8061
rect 3133 -8792 3199 -8782
rect 3325 -8071 3391 -8061
rect 3325 -8792 3391 -8782
rect 3517 -8071 3583 -8061
rect 3517 -8792 3583 -8782
rect 3709 -8071 3775 -8061
rect 3709 -8792 3775 -8782
rect 3901 -8071 3967 -8061
rect 3901 -8792 3967 -8782
rect 4093 -8071 4159 -8061
rect 4093 -8792 4159 -8782
rect 4285 -8071 4351 -8061
rect 4285 -8792 4351 -8782
rect 4477 -8071 4543 -8061
rect 4477 -8792 4543 -8782
rect 4669 -8071 4735 -8061
rect 4669 -8792 4735 -8782
rect 4861 -8071 4927 -8061
rect 4861 -8792 4927 -8782
rect 5053 -8071 5119 -8061
rect 5053 -8792 5119 -8782
rect 5245 -8071 5311 -8061
rect 5245 -8792 5311 -8782
rect 5437 -8071 5503 -8061
rect 5437 -8792 5503 -8782
rect 5691 -9007 5897 -7875
rect 6208 -8071 6414 -6564
rect 6198 -8782 6208 -8071
rect 6414 -8782 6424 -8071
rect -4375 -9071 -4149 -9007
rect -4375 -9181 -4365 -9071
rect -4159 -9181 -4149 -9071
rect -3933 -9073 -3923 -9017
rect -3857 -9073 -3847 -9017
rect -3741 -9073 -3731 -9017
rect -3665 -9073 -3655 -9017
rect -3549 -9073 -3539 -9017
rect -3473 -9073 -3463 -9017
rect -3357 -9073 -3347 -9017
rect -3281 -9073 -3271 -9017
rect -3165 -9073 -3155 -9017
rect -3089 -9073 -3079 -9017
rect -2973 -9073 -2963 -9017
rect -2897 -9073 -2887 -9017
rect -2781 -9073 -2771 -9017
rect -2705 -9073 -2695 -9017
rect -2589 -9073 -2579 -9017
rect -2513 -9073 -2503 -9017
rect -2397 -9073 -2387 -9017
rect -2321 -9073 -2311 -9017
rect -2205 -9073 -2195 -9017
rect -2129 -9073 -2119 -9017
rect -2013 -9073 -2003 -9017
rect -1937 -9073 -1927 -9017
rect -1821 -9073 -1811 -9017
rect -1745 -9073 -1735 -9017
rect -1629 -9073 -1619 -9017
rect -1553 -9073 -1543 -9017
rect -1437 -9073 -1427 -9017
rect -1361 -9073 -1351 -9017
rect -1245 -9073 -1235 -9017
rect -1169 -9073 -1159 -9017
rect -1053 -9073 -1043 -9017
rect -977 -9073 -967 -9017
rect -861 -9073 -851 -9017
rect -785 -9073 -775 -9017
rect -669 -9073 -659 -9017
rect -593 -9073 -583 -9017
rect -477 -9073 -467 -9017
rect -401 -9073 -391 -9017
rect -285 -9073 -275 -9017
rect -209 -9073 -199 -9017
rect -93 -9073 -83 -9017
rect -17 -9073 -7 -9017
rect 99 -9073 109 -9017
rect 175 -9073 185 -9017
rect 291 -9073 301 -9017
rect 367 -9073 377 -9017
rect 483 -9073 493 -9017
rect 559 -9073 569 -9017
rect 675 -9073 685 -9017
rect 751 -9073 761 -9017
rect 867 -9073 877 -9017
rect 943 -9073 953 -9017
rect 1059 -9073 1069 -9017
rect 1135 -9073 1145 -9017
rect 1251 -9073 1261 -9017
rect 1327 -9073 1337 -9017
rect 1443 -9073 1453 -9017
rect 1519 -9073 1529 -9017
rect 1635 -9073 1645 -9017
rect 1711 -9073 1721 -9017
rect 1827 -9073 1837 -9017
rect 1903 -9073 1913 -9017
rect 2019 -9073 2029 -9017
rect 2095 -9073 2105 -9017
rect 2211 -9073 2221 -9017
rect 2287 -9073 2297 -9017
rect 2403 -9073 2413 -9017
rect 2479 -9073 2489 -9017
rect 2595 -9073 2605 -9017
rect 2671 -9073 2681 -9017
rect 2787 -9073 2797 -9017
rect 2863 -9073 2873 -9017
rect 2979 -9073 2989 -9017
rect 3055 -9073 3065 -9017
rect 3171 -9073 3181 -9017
rect 3247 -9073 3257 -9017
rect 3363 -9073 3373 -9017
rect 3439 -9073 3449 -9017
rect 3555 -9073 3565 -9017
rect 3631 -9073 3641 -9017
rect 3747 -9073 3757 -9017
rect 3823 -9073 3833 -9017
rect 3939 -9073 3949 -9017
rect 4015 -9073 4025 -9017
rect 4131 -9073 4141 -9017
rect 4207 -9073 4217 -9017
rect 4323 -9073 4333 -9017
rect 4399 -9073 4409 -9017
rect 4515 -9073 4525 -9017
rect 4591 -9073 4601 -9017
rect 4707 -9073 4717 -9017
rect 4783 -9073 4793 -9017
rect 4899 -9073 4909 -9017
rect 4975 -9073 4985 -9017
rect 5091 -9073 5101 -9017
rect 5167 -9073 5177 -9017
rect 5283 -9073 5293 -9017
rect 5359 -9073 5369 -9017
rect 5475 -9073 5485 -9017
rect 5551 -9073 5561 -9017
rect -3933 -9171 -3923 -9115
rect -3857 -9171 -3847 -9115
rect -3741 -9171 -3731 -9115
rect -3665 -9171 -3655 -9115
rect -3549 -9171 -3539 -9115
rect -3473 -9171 -3463 -9115
rect -3357 -9171 -3347 -9115
rect -3281 -9171 -3271 -9115
rect -3165 -9171 -3155 -9115
rect -3089 -9171 -3079 -9115
rect -2973 -9171 -2963 -9115
rect -2897 -9171 -2887 -9115
rect -2781 -9171 -2771 -9115
rect -2705 -9171 -2695 -9115
rect -2589 -9171 -2579 -9115
rect -2513 -9171 -2503 -9115
rect -2397 -9171 -2387 -9115
rect -2321 -9171 -2311 -9115
rect -2205 -9171 -2195 -9115
rect -2129 -9171 -2119 -9115
rect -2013 -9171 -2003 -9115
rect -1937 -9171 -1927 -9115
rect -1821 -9171 -1811 -9115
rect -1745 -9171 -1735 -9115
rect -1629 -9171 -1619 -9115
rect -1553 -9171 -1543 -9115
rect -1437 -9171 -1427 -9115
rect -1361 -9171 -1351 -9115
rect -1245 -9171 -1235 -9115
rect -1169 -9171 -1159 -9115
rect -1053 -9171 -1043 -9115
rect -977 -9171 -967 -9115
rect -861 -9171 -851 -9115
rect -785 -9171 -775 -9115
rect -669 -9171 -659 -9115
rect -593 -9171 -583 -9115
rect -477 -9171 -467 -9115
rect -401 -9171 -391 -9115
rect -285 -9171 -275 -9115
rect -209 -9171 -199 -9115
rect -93 -9171 -83 -9115
rect -17 -9171 -7 -9115
rect 99 -9171 109 -9115
rect 175 -9171 185 -9115
rect 291 -9171 301 -9115
rect 367 -9171 377 -9115
rect 483 -9171 493 -9115
rect 559 -9171 569 -9115
rect 675 -9171 685 -9115
rect 751 -9171 761 -9115
rect 867 -9171 877 -9115
rect 943 -9171 953 -9115
rect 1059 -9171 1069 -9115
rect 1135 -9171 1145 -9115
rect 1251 -9171 1261 -9115
rect 1327 -9171 1337 -9115
rect 1443 -9171 1453 -9115
rect 1519 -9171 1529 -9115
rect 1635 -9171 1645 -9115
rect 1711 -9171 1721 -9115
rect 1827 -9171 1837 -9115
rect 1903 -9171 1913 -9115
rect 2019 -9171 2029 -9115
rect 2095 -9171 2105 -9115
rect 2211 -9171 2221 -9115
rect 2287 -9171 2297 -9115
rect 2403 -9171 2413 -9115
rect 2479 -9171 2489 -9115
rect 2595 -9171 2605 -9115
rect 2671 -9171 2681 -9115
rect 2787 -9171 2797 -9115
rect 2863 -9171 2873 -9115
rect 2979 -9171 2989 -9115
rect 3055 -9171 3065 -9115
rect 3171 -9171 3181 -9115
rect 3247 -9171 3257 -9115
rect 3363 -9171 3373 -9115
rect 3439 -9171 3449 -9115
rect 3555 -9171 3565 -9115
rect 3631 -9171 3641 -9115
rect 3747 -9171 3757 -9115
rect 3823 -9171 3833 -9115
rect 3939 -9171 3949 -9115
rect 4015 -9171 4025 -9115
rect 4131 -9171 4141 -9115
rect 4207 -9171 4217 -9115
rect 4323 -9171 4333 -9115
rect 4399 -9171 4409 -9115
rect 4515 -9171 4525 -9115
rect 4591 -9171 4601 -9115
rect 4707 -9171 4717 -9115
rect 4783 -9171 4793 -9115
rect 4899 -9171 4909 -9115
rect 4975 -9171 4985 -9115
rect 5091 -9171 5101 -9115
rect 5167 -9171 5177 -9115
rect 5283 -9171 5293 -9115
rect 5359 -9171 5369 -9115
rect 5475 -9171 5485 -9115
rect 5551 -9171 5561 -9115
rect 5681 -9181 5691 -9007
rect 5897 -9181 5907 -9007
rect -4365 -9392 -4159 -9181
rect -4063 -9392 -4011 -9382
rect -4375 -10093 -4365 -9392
rect -4159 -10093 -4149 -9392
rect -4800 -11000 -4790 -10289
rect -4584 -11000 -4574 -10289
rect -4791 -11399 -4584 -11000
rect -4365 -11225 -4159 -10093
rect -4063 -10103 -4011 -10093
rect -3871 -9392 -3819 -9382
rect -3871 -10103 -3819 -10093
rect -3679 -9392 -3627 -9382
rect -3679 -10103 -3627 -10093
rect -3487 -9392 -3435 -9382
rect -3487 -10103 -3435 -10093
rect -3295 -9392 -3243 -9382
rect -3295 -10103 -3243 -10093
rect -3103 -9392 -3051 -9382
rect -3103 -10103 -3051 -10093
rect -2911 -9392 -2859 -9382
rect -2911 -10103 -2859 -10093
rect -2719 -9392 -2667 -9382
rect -2719 -10103 -2667 -10093
rect -2527 -9392 -2475 -9382
rect -2527 -10103 -2475 -10093
rect -2335 -9392 -2283 -9382
rect -2335 -10103 -2283 -10093
rect -2143 -9392 -2091 -9382
rect -2143 -10103 -2091 -10093
rect -1951 -9392 -1899 -9382
rect -1951 -10103 -1899 -10093
rect -1759 -9392 -1707 -9382
rect -1759 -10103 -1707 -10093
rect -1567 -9392 -1515 -9382
rect -1567 -10103 -1515 -10093
rect -1375 -9392 -1323 -9382
rect -1375 -10103 -1323 -10093
rect -1183 -9392 -1131 -9382
rect -1183 -10103 -1131 -10093
rect -991 -9392 -939 -9382
rect -991 -10103 -939 -10093
rect -799 -9392 -747 -9382
rect -799 -10103 -747 -10093
rect -607 -9392 -555 -9382
rect -607 -10103 -555 -10093
rect -415 -9392 -363 -9382
rect -415 -10103 -363 -10093
rect -223 -9392 -171 -9382
rect -223 -10103 -171 -10093
rect -31 -9392 21 -9382
rect -31 -10103 21 -10093
rect 161 -9392 213 -9382
rect 161 -10103 213 -10093
rect 353 -9392 405 -9382
rect 353 -10103 405 -10093
rect 545 -9392 597 -9382
rect 545 -10103 597 -10093
rect 737 -9392 789 -9382
rect 737 -10103 789 -10093
rect 929 -9392 981 -9382
rect 929 -10103 981 -10093
rect 1121 -9392 1173 -9382
rect 1121 -10103 1173 -10093
rect 1313 -9392 1365 -9382
rect 1313 -10103 1365 -10093
rect 1505 -9392 1557 -9382
rect 1505 -10103 1557 -10093
rect 1697 -9392 1749 -9382
rect 1697 -10103 1749 -10093
rect 1889 -9392 1941 -9382
rect 1889 -10103 1941 -10093
rect 2081 -9392 2133 -9382
rect 2081 -10103 2133 -10093
rect 2273 -9392 2325 -9382
rect 2273 -10103 2325 -10093
rect 2465 -9392 2517 -9382
rect 2465 -10103 2517 -10093
rect 2657 -9392 2709 -9382
rect 2657 -10103 2709 -10093
rect 2849 -9392 2901 -9382
rect 2849 -10103 2901 -10093
rect 3041 -9392 3093 -9382
rect 3041 -10103 3093 -10093
rect 3233 -9392 3285 -9382
rect 3233 -10103 3285 -10093
rect 3425 -9392 3477 -9382
rect 3425 -10103 3477 -10093
rect 3617 -9392 3669 -9382
rect 3617 -10103 3669 -10093
rect 3809 -9392 3861 -9382
rect 3809 -10103 3861 -10093
rect 4001 -9392 4053 -9382
rect 4001 -10103 4053 -10093
rect 4193 -9392 4245 -9382
rect 4193 -10103 4245 -10093
rect 4385 -9392 4437 -9382
rect 4385 -10103 4437 -10093
rect 4577 -9392 4629 -9382
rect 4577 -10103 4629 -10093
rect 4769 -9392 4821 -9382
rect 4769 -10103 4821 -10093
rect 4961 -9392 5013 -9382
rect 4961 -10103 5013 -10093
rect 5153 -9392 5205 -9382
rect 5153 -10103 5205 -10093
rect 5345 -9392 5397 -9382
rect 5691 -9392 5897 -9181
rect 5527 -10093 5537 -9392
rect 5589 -10093 5599 -9392
rect 5681 -10093 5691 -9392
rect 5897 -10093 5907 -9392
rect 5345 -10103 5397 -10093
rect -3971 -10289 -3905 -10279
rect -3971 -11010 -3905 -11000
rect -3779 -10289 -3713 -10279
rect -3779 -11010 -3713 -11000
rect -3587 -10289 -3521 -10279
rect -3587 -11010 -3521 -11000
rect -3395 -10289 -3329 -10279
rect -3395 -11010 -3329 -11000
rect -3203 -10289 -3137 -10279
rect -3203 -11010 -3137 -11000
rect -3011 -10289 -2945 -10279
rect -3011 -11010 -2945 -11000
rect -2819 -10289 -2753 -10279
rect -2819 -11010 -2753 -11000
rect -2627 -10289 -2561 -10279
rect -2627 -11010 -2561 -11000
rect -2435 -10289 -2369 -10279
rect -2435 -11010 -2369 -11000
rect -2243 -10289 -2177 -10279
rect -2243 -11010 -2177 -11000
rect -2051 -10289 -1985 -10279
rect -2051 -11010 -1985 -11000
rect -1859 -10289 -1793 -10279
rect -1859 -11010 -1793 -11000
rect -1667 -10289 -1601 -10279
rect -1667 -11010 -1601 -11000
rect -1475 -10289 -1409 -10279
rect -1475 -11010 -1409 -11000
rect -1283 -10289 -1217 -10279
rect -1283 -11010 -1217 -11000
rect -1091 -10289 -1025 -10279
rect -1091 -11010 -1025 -11000
rect -899 -10289 -833 -10279
rect -899 -11010 -833 -11000
rect -707 -10289 -641 -10279
rect -707 -11010 -641 -11000
rect -515 -10289 -449 -10279
rect -515 -11010 -449 -11000
rect -323 -10289 -257 -10279
rect -323 -11010 -257 -11000
rect -131 -10289 -65 -10279
rect -131 -11010 -65 -11000
rect 61 -10289 127 -10279
rect 61 -11010 127 -11000
rect 253 -10289 319 -10279
rect 253 -11010 319 -11000
rect 445 -10289 511 -10279
rect 445 -11010 511 -11000
rect 637 -10289 703 -10279
rect 637 -11010 703 -11000
rect 829 -10289 895 -10279
rect 829 -11010 895 -11000
rect 1021 -10289 1087 -10279
rect 1021 -11010 1087 -11000
rect 1213 -10289 1279 -10279
rect 1213 -11010 1279 -11000
rect 1405 -10289 1471 -10279
rect 1405 -11010 1471 -11000
rect 1597 -10289 1663 -10279
rect 1597 -11010 1663 -11000
rect 1789 -10289 1855 -10279
rect 1789 -11010 1855 -11000
rect 1981 -10289 2047 -10279
rect 1981 -11010 2047 -11000
rect 2173 -10289 2239 -10279
rect 2173 -11010 2239 -11000
rect 2365 -10289 2431 -10279
rect 2365 -11010 2431 -11000
rect 2557 -10289 2623 -10279
rect 2557 -11010 2623 -11000
rect 2749 -10289 2815 -10279
rect 2749 -11010 2815 -11000
rect 2941 -10289 3007 -10279
rect 2941 -11010 3007 -11000
rect 3133 -10289 3199 -10279
rect 3133 -11010 3199 -11000
rect 3325 -10289 3391 -10279
rect 3325 -11010 3391 -11000
rect 3517 -10289 3583 -10279
rect 3517 -11010 3583 -11000
rect 3709 -10289 3775 -10279
rect 3709 -11010 3775 -11000
rect 3901 -10289 3967 -10279
rect 3901 -11010 3967 -11000
rect 4093 -10289 4159 -10279
rect 4093 -11010 4159 -11000
rect 4285 -10289 4351 -10279
rect 4285 -11010 4351 -11000
rect 4477 -10289 4543 -10279
rect 4477 -11010 4543 -11000
rect 4669 -10289 4735 -10279
rect 4669 -11010 4735 -11000
rect 4861 -10289 4927 -10279
rect 4861 -11010 4927 -11000
rect 5053 -10289 5119 -10279
rect 5053 -11010 5119 -11000
rect 5245 -10289 5311 -10279
rect 5245 -11010 5311 -11000
rect 5437 -10289 5503 -10279
rect 5437 -11010 5503 -11000
rect 5691 -11225 5897 -10093
rect 6208 -10289 6414 -8782
rect 6198 -11000 6208 -10289
rect 6414 -11000 6424 -10289
rect -4375 -11399 -4365 -11225
rect -4159 -11399 -4149 -11225
rect -4029 -11291 -4019 -11235
rect -3953 -11291 -3943 -11235
rect -3837 -11291 -3827 -11235
rect -3761 -11291 -3751 -11235
rect -3645 -11291 -3635 -11235
rect -3569 -11291 -3559 -11235
rect -3453 -11291 -3443 -11235
rect -3377 -11291 -3367 -11235
rect -3261 -11291 -3251 -11235
rect -3185 -11291 -3175 -11235
rect -3069 -11291 -3059 -11235
rect -2993 -11291 -2983 -11235
rect -2877 -11291 -2867 -11235
rect -2801 -11291 -2791 -11235
rect -2685 -11291 -2675 -11235
rect -2609 -11291 -2599 -11235
rect -2493 -11291 -2483 -11235
rect -2417 -11291 -2407 -11235
rect -2301 -11291 -2291 -11235
rect -2225 -11291 -2215 -11235
rect -2109 -11291 -2099 -11235
rect -2033 -11291 -2023 -11235
rect -1917 -11291 -1907 -11235
rect -1841 -11291 -1831 -11235
rect -1725 -11291 -1715 -11235
rect -1649 -11291 -1639 -11235
rect -1533 -11291 -1523 -11235
rect -1457 -11291 -1447 -11235
rect -1341 -11291 -1331 -11235
rect -1265 -11291 -1255 -11235
rect -1149 -11291 -1139 -11235
rect -1073 -11291 -1063 -11235
rect -957 -11291 -947 -11235
rect -881 -11291 -871 -11235
rect -765 -11291 -755 -11235
rect -689 -11291 -679 -11235
rect -573 -11291 -563 -11235
rect -497 -11291 -487 -11235
rect -381 -11291 -371 -11235
rect -305 -11291 -295 -11235
rect -189 -11291 -179 -11235
rect -113 -11291 -103 -11235
rect 3 -11291 13 -11235
rect 79 -11291 89 -11235
rect 195 -11291 205 -11235
rect 271 -11291 281 -11235
rect 387 -11291 397 -11235
rect 463 -11291 473 -11235
rect 579 -11291 589 -11235
rect 655 -11291 665 -11235
rect 771 -11291 781 -11235
rect 847 -11291 857 -11235
rect 963 -11291 973 -11235
rect 1039 -11291 1049 -11235
rect 1155 -11291 1165 -11235
rect 1231 -11291 1241 -11235
rect 1347 -11291 1357 -11235
rect 1423 -11291 1433 -11235
rect 1539 -11291 1549 -11235
rect 1615 -11291 1625 -11235
rect 1731 -11291 1741 -11235
rect 1807 -11291 1817 -11235
rect 1923 -11291 1933 -11235
rect 1999 -11291 2009 -11235
rect 2115 -11291 2125 -11235
rect 2191 -11291 2201 -11235
rect 2307 -11291 2317 -11235
rect 2383 -11291 2393 -11235
rect 2499 -11291 2509 -11235
rect 2575 -11291 2585 -11235
rect 2691 -11291 2701 -11235
rect 2767 -11291 2777 -11235
rect 2883 -11291 2893 -11235
rect 2959 -11291 2969 -11235
rect 3075 -11291 3085 -11235
rect 3151 -11291 3161 -11235
rect 3267 -11291 3277 -11235
rect 3343 -11291 3353 -11235
rect 3459 -11291 3469 -11235
rect 3535 -11291 3545 -11235
rect 3651 -11291 3661 -11235
rect 3727 -11291 3737 -11235
rect 3843 -11291 3853 -11235
rect 3919 -11291 3929 -11235
rect 4035 -11291 4045 -11235
rect 4111 -11291 4121 -11235
rect 4227 -11291 4237 -11235
rect 4303 -11291 4313 -11235
rect 4419 -11291 4429 -11235
rect 4495 -11291 4505 -11235
rect 4611 -11291 4621 -11235
rect 4687 -11291 4697 -11235
rect 4803 -11291 4813 -11235
rect 4879 -11291 4889 -11235
rect 4995 -11291 5005 -11235
rect 5071 -11291 5081 -11235
rect 5187 -11291 5197 -11235
rect 5263 -11291 5273 -11235
rect 5379 -11291 5389 -11235
rect 5455 -11291 5465 -11235
rect 5681 -11399 5691 -11225
rect 5897 -11399 5907 -11225
rect 6208 -11399 6414 -11000
<< via1 >>
rect -3193 1076 -2900 1369
rect 29 1066 87 1366
rect 383 1435 441 1715
rect 265 1066 323 1366
rect 147 715 205 1015
rect 501 1066 559 1366
rect 855 1435 913 1715
rect 737 1066 795 1366
rect 619 715 677 1015
rect 973 1066 1031 1366
rect 1327 1435 1385 1715
rect 1209 1066 1267 1366
rect 1091 715 1149 1015
rect 1445 1066 1503 1366
rect 4442 1076 4735 1369
rect 321 69 1211 225
rect -2678 -268 -2619 -202
rect -823 -268 -764 -202
rect -2222 -599 -2164 -299
rect -1750 -599 -1692 -299
rect -1278 -599 -1220 -299
rect -2678 -949 -2619 -649
rect -2458 -949 -2400 -649
rect -1986 -949 -1928 -649
rect -1514 -949 -1456 -649
rect -1042 -949 -984 -649
rect -823 -949 -764 -649
rect -2576 -1299 -2518 -999
rect -2340 -1299 -2282 -999
rect -2104 -1299 -2046 -999
rect -1868 -1299 -1810 -999
rect -1632 -1299 -1574 -999
rect -1396 -1299 -1338 -999
rect -1160 -1299 -1102 -999
rect -924 -1299 -866 -999
rect -2678 -1396 -2619 -1337
rect -2403 -1396 -1039 -1337
rect -53 -1090 5 -527
rect -823 -1396 -764 -1337
rect 105 -1599 163 -1145
rect 263 -1090 321 -527
rect 421 -472 479 -18
rect 579 -1090 637 -527
rect 895 -1090 953 -527
rect 737 -1599 795 -1145
rect 1053 -472 1111 -18
rect 1211 -1090 1269 -527
rect 1369 -1599 1427 -1145
rect 2296 -268 2355 -202
rect 1527 -1090 1585 -527
rect 4151 -268 4210 -202
rect 2752 -599 2810 -299
rect 3224 -599 3282 -299
rect 3696 -599 3754 -299
rect 2296 -949 2355 -649
rect 2516 -949 2574 -649
rect 2988 -949 3046 -649
rect 3460 -949 3518 -649
rect 3932 -949 3990 -649
rect 4151 -949 4210 -649
rect 2398 -1299 2456 -999
rect 2634 -1299 2692 -999
rect 2870 -1299 2928 -999
rect 3106 -1299 3164 -999
rect 3342 -1299 3400 -999
rect 3578 -1299 3636 -999
rect 3814 -1299 3872 -999
rect 4050 -1299 4108 -999
rect 2296 -1396 2355 -1337
rect 2571 -1396 3935 -1337
rect 4151 -1396 4210 -1337
rect 163 -1823 1369 -1667
rect -1932 -2597 -1707 -2382
rect -1259 -2394 2791 -2382
rect -1259 -2537 -1247 -2394
rect -1247 -2537 2779 -2394
rect 2779 -2537 2791 -2394
rect -1259 -2607 2791 -2537
rect 3249 -2603 3474 -2388
rect -1327 -2948 -1269 -2655
rect -295 -2948 -237 -2655
rect 737 -2948 795 -2655
rect 1769 -2948 1827 -2655
rect 2801 -2948 2859 -2655
rect -1932 -3294 -1707 -2996
rect -811 -3294 -753 -2996
rect 221 -3294 279 -2996
rect 1253 -3294 1311 -2996
rect 2285 -3294 2343 -2996
rect 3249 -3294 3474 -2996
rect -3193 -3635 -2900 -3342
rect -2091 -3645 -2041 -3332
rect -2041 -3645 -2007 -3332
rect -2007 -3645 -2001 -3332
rect -1585 -3635 -1527 -3342
rect -1069 -3635 -1011 -3342
rect -553 -3635 -495 -3342
rect -37 -3635 21 -3342
rect 479 -3635 537 -3342
rect 995 -3635 1053 -3342
rect 1511 -3635 1569 -3342
rect 2027 -3635 2085 -3342
rect 2543 -3635 2601 -3342
rect 3059 -3635 3117 -3342
rect -1932 -3908 -1707 -3683
rect -1259 -3753 2791 -3683
rect -1259 -3896 -1247 -3753
rect -1247 -3896 2779 -3753
rect 2779 -3896 2791 -3753
rect -1259 -3908 2791 -3896
rect 3543 -3645 3549 -3332
rect 3549 -3645 3583 -3332
rect 3583 -3645 3633 -3332
rect 4442 -3635 4735 -3342
rect 3249 -3908 3474 -3693
rect -4791 -4435 -4584 -4262
rect 6208 -4435 6415 -4262
rect -4974 -5657 -4940 -4571
rect -4940 -5657 -4875 -4571
rect -4875 -5657 -4841 -4571
rect -4365 -4745 -4159 -4571
rect -3923 -4735 -3857 -4679
rect -3731 -4735 -3665 -4679
rect -3539 -4735 -3473 -4679
rect -3347 -4735 -3281 -4679
rect -3155 -4735 -3089 -4679
rect -2963 -4735 -2897 -4679
rect -2771 -4735 -2705 -4679
rect -2579 -4735 -2513 -4679
rect -2387 -4735 -2321 -4679
rect -2195 -4735 -2129 -4679
rect -2003 -4735 -1937 -4679
rect -1811 -4735 -1745 -4679
rect -1619 -4735 -1553 -4679
rect -1427 -4735 -1361 -4679
rect -1235 -4735 -1169 -4679
rect -1043 -4735 -977 -4679
rect -851 -4735 -785 -4679
rect -659 -4735 -593 -4679
rect -467 -4735 -401 -4679
rect -275 -4735 -209 -4679
rect -83 -4735 -17 -4679
rect 109 -4735 175 -4679
rect 301 -4735 367 -4679
rect 493 -4735 559 -4679
rect 685 -4735 751 -4679
rect 877 -4735 943 -4679
rect 1069 -4735 1135 -4679
rect 1261 -4735 1327 -4679
rect 1453 -4735 1519 -4679
rect 1645 -4735 1711 -4679
rect 1837 -4735 1903 -4679
rect 2029 -4735 2095 -4679
rect 2221 -4735 2287 -4679
rect 2413 -4735 2479 -4679
rect 2605 -4735 2671 -4679
rect 2797 -4735 2863 -4679
rect 2989 -4735 3055 -4679
rect 3181 -4735 3247 -4679
rect 3373 -4735 3439 -4679
rect 3565 -4735 3631 -4679
rect 3757 -4735 3823 -4679
rect 3949 -4735 4015 -4679
rect 4141 -4735 4207 -4679
rect 4333 -4735 4399 -4679
rect 4525 -4735 4591 -4679
rect 4717 -4735 4783 -4679
rect 4909 -4735 4975 -4679
rect 5101 -4735 5167 -4679
rect 5293 -4735 5359 -4679
rect 5485 -4735 5551 -4679
rect 5691 -4745 5897 -4571
rect -4365 -5657 -4159 -4956
rect -4063 -5657 -4011 -4956
rect -4790 -6564 -4584 -5853
rect -3871 -5657 -3819 -4956
rect -3679 -5657 -3627 -4956
rect -3487 -5657 -3435 -4956
rect -3295 -5657 -3243 -4956
rect -3103 -5657 -3051 -4956
rect -2911 -5657 -2859 -4956
rect -2719 -5657 -2667 -4956
rect -2527 -5657 -2475 -4956
rect -2335 -5657 -2283 -4956
rect -2143 -5657 -2091 -4956
rect -1951 -5657 -1899 -4956
rect -1759 -5657 -1707 -4956
rect -1567 -5657 -1515 -4956
rect -1375 -5657 -1323 -4956
rect -1183 -5657 -1131 -4956
rect -991 -5657 -939 -4956
rect -799 -5657 -747 -4956
rect -607 -5657 -555 -4956
rect -415 -5657 -363 -4956
rect -223 -5657 -171 -4956
rect -31 -5657 21 -4956
rect 161 -5657 213 -4956
rect 353 -5657 405 -4956
rect 545 -5657 597 -4956
rect 737 -5657 789 -4956
rect 929 -5657 981 -4956
rect 1121 -5657 1173 -4956
rect 1313 -5657 1365 -4956
rect 1505 -5657 1557 -4956
rect 1697 -5657 1749 -4956
rect 1889 -5657 1941 -4956
rect 2081 -5657 2133 -4956
rect 2273 -5657 2325 -4956
rect 2465 -5657 2517 -4956
rect 2657 -5657 2709 -4956
rect 2849 -5657 2901 -4956
rect 3041 -5657 3093 -4956
rect 3233 -5657 3285 -4956
rect 3425 -5657 3477 -4956
rect 3617 -5657 3669 -4956
rect 3809 -5657 3861 -4956
rect 4001 -5657 4053 -4956
rect 4193 -5657 4245 -4956
rect 4385 -5657 4437 -4956
rect 4577 -5657 4629 -4956
rect 4769 -5657 4821 -4956
rect 4961 -5657 5013 -4956
rect 5153 -5657 5205 -4956
rect 5345 -5657 5397 -4956
rect 5537 -5657 5589 -4956
rect 5691 -5657 5897 -4956
rect -3971 -6564 -3905 -5853
rect -3779 -6564 -3713 -5853
rect -3587 -6564 -3521 -5853
rect -3395 -6564 -3329 -5853
rect -3203 -6564 -3137 -5853
rect -3011 -6564 -2945 -5853
rect -2819 -6564 -2753 -5853
rect -2627 -6564 -2561 -5853
rect -2435 -6564 -2369 -5853
rect -2243 -6564 -2177 -5853
rect -2051 -6564 -1985 -5853
rect -1859 -6564 -1793 -5853
rect -1667 -6564 -1601 -5853
rect -1475 -6564 -1409 -5853
rect -1283 -6564 -1217 -5853
rect -1091 -6564 -1025 -5853
rect -899 -6564 -833 -5853
rect -707 -6564 -641 -5853
rect -515 -6564 -449 -5853
rect -323 -6564 -257 -5853
rect -131 -6564 -65 -5853
rect 61 -6564 127 -5853
rect 253 -6564 319 -5853
rect 445 -6564 511 -5853
rect 637 -6564 703 -5853
rect 829 -6564 895 -5853
rect 1021 -6564 1087 -5853
rect 1213 -6564 1279 -5853
rect 1405 -6564 1471 -5853
rect 1597 -6564 1663 -5853
rect 1789 -6564 1855 -5853
rect 1981 -6564 2047 -5853
rect 2173 -6564 2239 -5853
rect 2365 -6564 2431 -5853
rect 2557 -6564 2623 -5853
rect 2749 -6564 2815 -5853
rect 2941 -6564 3007 -5853
rect 3133 -6564 3199 -5853
rect 3325 -6564 3391 -5853
rect 3517 -6564 3583 -5853
rect 3709 -6564 3775 -5853
rect 3901 -6564 3967 -5853
rect 4093 -6564 4159 -5853
rect 4285 -6564 4351 -5853
rect 4477 -6564 4543 -5853
rect 4669 -6564 4735 -5853
rect 4861 -6564 4927 -5853
rect 5053 -6564 5119 -5853
rect 5245 -6564 5311 -5853
rect 5437 -6564 5503 -5853
rect 6465 -5657 6499 -4571
rect 6499 -5657 6563 -4571
rect 6563 -5657 6597 -4571
rect 6597 -5657 6598 -4571
rect 6208 -6564 6414 -5853
rect -4365 -6963 -4159 -6789
rect -4019 -6855 -3953 -6799
rect -3827 -6855 -3761 -6799
rect -3635 -6855 -3569 -6799
rect -3443 -6855 -3377 -6799
rect -3251 -6855 -3185 -6799
rect -3059 -6855 -2993 -6799
rect -2867 -6855 -2801 -6799
rect -2675 -6855 -2609 -6799
rect -2483 -6855 -2417 -6799
rect -2291 -6855 -2225 -6799
rect -2099 -6855 -2033 -6799
rect -1907 -6855 -1841 -6799
rect -1715 -6855 -1649 -6799
rect -1523 -6855 -1457 -6799
rect -1331 -6855 -1265 -6799
rect -1139 -6855 -1073 -6799
rect -947 -6855 -881 -6799
rect -755 -6855 -689 -6799
rect -563 -6855 -497 -6799
rect -371 -6855 -305 -6799
rect -179 -6855 -113 -6799
rect 13 -6855 79 -6799
rect 205 -6855 271 -6799
rect 397 -6855 463 -6799
rect 589 -6855 655 -6799
rect 781 -6855 847 -6799
rect 973 -6855 1039 -6799
rect 1165 -6855 1231 -6799
rect 1357 -6855 1423 -6799
rect 1549 -6855 1615 -6799
rect 1741 -6855 1807 -6799
rect 1933 -6855 1999 -6799
rect 2125 -6855 2191 -6799
rect 2317 -6855 2383 -6799
rect 2509 -6855 2575 -6799
rect 2701 -6855 2767 -6799
rect 2893 -6855 2959 -6799
rect 3085 -6855 3151 -6799
rect 3277 -6855 3343 -6799
rect 3469 -6855 3535 -6799
rect 3661 -6855 3727 -6799
rect 3853 -6855 3919 -6799
rect 4045 -6855 4111 -6799
rect 4237 -6855 4303 -6799
rect 4429 -6855 4495 -6799
rect 4621 -6855 4687 -6799
rect 4813 -6855 4879 -6799
rect 5005 -6855 5071 -6799
rect 5197 -6855 5263 -6799
rect 5389 -6855 5455 -6799
rect -4019 -6953 -3953 -6897
rect -3827 -6953 -3761 -6897
rect -3635 -6953 -3569 -6897
rect -3443 -6953 -3377 -6897
rect -3251 -6953 -3185 -6897
rect -3059 -6953 -2993 -6897
rect -2867 -6953 -2801 -6897
rect -2675 -6953 -2609 -6897
rect -2483 -6953 -2417 -6897
rect -2291 -6953 -2225 -6897
rect -2099 -6953 -2033 -6897
rect -1907 -6953 -1841 -6897
rect -1715 -6953 -1649 -6897
rect -1523 -6953 -1457 -6897
rect -1331 -6953 -1265 -6897
rect -1139 -6953 -1073 -6897
rect -947 -6953 -881 -6897
rect -755 -6953 -689 -6897
rect -563 -6953 -497 -6897
rect -371 -6953 -305 -6897
rect -179 -6953 -113 -6897
rect 13 -6953 79 -6897
rect 205 -6953 271 -6897
rect 397 -6953 463 -6897
rect 589 -6953 655 -6897
rect 781 -6953 847 -6897
rect 973 -6953 1039 -6897
rect 1165 -6953 1231 -6897
rect 1357 -6953 1423 -6897
rect 1549 -6953 1615 -6897
rect 1741 -6953 1807 -6897
rect 1933 -6953 1999 -6897
rect 2125 -6953 2191 -6897
rect 2317 -6953 2383 -6897
rect 2509 -6953 2575 -6897
rect 2701 -6953 2767 -6897
rect 2893 -6953 2959 -6897
rect 3085 -6953 3151 -6897
rect 3277 -6953 3343 -6897
rect 3469 -6953 3535 -6897
rect 3661 -6953 3727 -6897
rect 3853 -6953 3919 -6897
rect 4045 -6953 4111 -6897
rect 4237 -6953 4303 -6897
rect 4429 -6953 4495 -6897
rect 4621 -6953 4687 -6897
rect 4813 -6953 4879 -6897
rect 5005 -6953 5071 -6897
rect 5197 -6953 5263 -6897
rect 5389 -6953 5455 -6897
rect 5691 -6963 5897 -6789
rect -4365 -7875 -4159 -7174
rect -4063 -7875 -4011 -7174
rect -4790 -8782 -4584 -8071
rect -3871 -7875 -3819 -7174
rect -3679 -7875 -3627 -7174
rect -3487 -7875 -3435 -7174
rect -3295 -7875 -3243 -7174
rect -3103 -7875 -3051 -7174
rect -2911 -7875 -2859 -7174
rect -2719 -7875 -2667 -7174
rect -2527 -7875 -2475 -7174
rect -2335 -7875 -2283 -7174
rect -2143 -7875 -2091 -7174
rect -1951 -7875 -1899 -7174
rect -1759 -7875 -1707 -7174
rect -1567 -7875 -1515 -7174
rect -1375 -7875 -1323 -7174
rect -1183 -7875 -1131 -7174
rect -991 -7875 -939 -7174
rect -799 -7875 -747 -7174
rect -607 -7875 -555 -7174
rect -415 -7875 -363 -7174
rect -223 -7875 -171 -7174
rect -31 -7875 21 -7174
rect 161 -7875 213 -7174
rect 353 -7875 405 -7174
rect 545 -7875 597 -7174
rect 737 -7875 789 -7174
rect 929 -7875 981 -7174
rect 1121 -7875 1173 -7174
rect 1313 -7875 1365 -7174
rect 1505 -7875 1557 -7174
rect 1697 -7875 1749 -7174
rect 1889 -7875 1941 -7174
rect 2081 -7875 2133 -7174
rect 2273 -7875 2325 -7174
rect 2465 -7875 2517 -7174
rect 2657 -7875 2709 -7174
rect 2849 -7875 2901 -7174
rect 3041 -7875 3093 -7174
rect 3233 -7875 3285 -7174
rect 3425 -7875 3477 -7174
rect 3617 -7875 3669 -7174
rect 3809 -7875 3861 -7174
rect 4001 -7875 4053 -7174
rect 4193 -7875 4245 -7174
rect 4385 -7875 4437 -7174
rect 4577 -7875 4629 -7174
rect 4769 -7875 4821 -7174
rect 4961 -7875 5013 -7174
rect 5153 -7875 5205 -7174
rect 5345 -7875 5397 -7174
rect 5537 -7875 5589 -7174
rect 5691 -7875 5897 -7174
rect -3971 -8782 -3905 -8071
rect -3779 -8782 -3713 -8071
rect -3587 -8782 -3521 -8071
rect -3395 -8782 -3329 -8071
rect -3203 -8782 -3137 -8071
rect -3011 -8782 -2945 -8071
rect -2819 -8782 -2753 -8071
rect -2627 -8782 -2561 -8071
rect -2435 -8782 -2369 -8071
rect -2243 -8782 -2177 -8071
rect -2051 -8782 -1985 -8071
rect -1859 -8782 -1793 -8071
rect -1667 -8782 -1601 -8071
rect -1475 -8782 -1409 -8071
rect -1283 -8782 -1217 -8071
rect -1091 -8782 -1025 -8071
rect -899 -8782 -833 -8071
rect -707 -8782 -641 -8071
rect -515 -8782 -449 -8071
rect -323 -8782 -257 -8071
rect -131 -8782 -65 -8071
rect 61 -8782 127 -8071
rect 253 -8782 319 -8071
rect 445 -8782 511 -8071
rect 637 -8782 703 -8071
rect 829 -8782 895 -8071
rect 1021 -8782 1087 -8071
rect 1213 -8782 1279 -8071
rect 1405 -8782 1471 -8071
rect 1597 -8782 1663 -8071
rect 1789 -8782 1855 -8071
rect 1981 -8782 2047 -8071
rect 2173 -8782 2239 -8071
rect 2365 -8782 2431 -8071
rect 2557 -8782 2623 -8071
rect 2749 -8782 2815 -8071
rect 2941 -8782 3007 -8071
rect 3133 -8782 3199 -8071
rect 3325 -8782 3391 -8071
rect 3517 -8782 3583 -8071
rect 3709 -8782 3775 -8071
rect 3901 -8782 3967 -8071
rect 4093 -8782 4159 -8071
rect 4285 -8782 4351 -8071
rect 4477 -8782 4543 -8071
rect 4669 -8782 4735 -8071
rect 4861 -8782 4927 -8071
rect 5053 -8782 5119 -8071
rect 5245 -8782 5311 -8071
rect 5437 -8782 5503 -8071
rect 6208 -8782 6414 -8071
rect -4365 -9181 -4159 -9071
rect -3923 -9073 -3857 -9017
rect -3731 -9073 -3665 -9017
rect -3539 -9073 -3473 -9017
rect -3347 -9073 -3281 -9017
rect -3155 -9073 -3089 -9017
rect -2963 -9073 -2897 -9017
rect -2771 -9073 -2705 -9017
rect -2579 -9073 -2513 -9017
rect -2387 -9073 -2321 -9017
rect -2195 -9073 -2129 -9017
rect -2003 -9073 -1937 -9017
rect -1811 -9073 -1745 -9017
rect -1619 -9073 -1553 -9017
rect -1427 -9073 -1361 -9017
rect -1235 -9073 -1169 -9017
rect -1043 -9073 -977 -9017
rect -851 -9073 -785 -9017
rect -659 -9073 -593 -9017
rect -467 -9073 -401 -9017
rect -275 -9073 -209 -9017
rect -83 -9073 -17 -9017
rect 109 -9073 175 -9017
rect 301 -9073 367 -9017
rect 493 -9073 559 -9017
rect 685 -9073 751 -9017
rect 877 -9073 943 -9017
rect 1069 -9073 1135 -9017
rect 1261 -9073 1327 -9017
rect 1453 -9073 1519 -9017
rect 1645 -9073 1711 -9017
rect 1837 -9073 1903 -9017
rect 2029 -9073 2095 -9017
rect 2221 -9073 2287 -9017
rect 2413 -9073 2479 -9017
rect 2605 -9073 2671 -9017
rect 2797 -9073 2863 -9017
rect 2989 -9073 3055 -9017
rect 3181 -9073 3247 -9017
rect 3373 -9073 3439 -9017
rect 3565 -9073 3631 -9017
rect 3757 -9073 3823 -9017
rect 3949 -9073 4015 -9017
rect 4141 -9073 4207 -9017
rect 4333 -9073 4399 -9017
rect 4525 -9073 4591 -9017
rect 4717 -9073 4783 -9017
rect 4909 -9073 4975 -9017
rect 5101 -9073 5167 -9017
rect 5293 -9073 5359 -9017
rect 5485 -9073 5551 -9017
rect -3923 -9171 -3857 -9115
rect -3731 -9171 -3665 -9115
rect -3539 -9171 -3473 -9115
rect -3347 -9171 -3281 -9115
rect -3155 -9171 -3089 -9115
rect -2963 -9171 -2897 -9115
rect -2771 -9171 -2705 -9115
rect -2579 -9171 -2513 -9115
rect -2387 -9171 -2321 -9115
rect -2195 -9171 -2129 -9115
rect -2003 -9171 -1937 -9115
rect -1811 -9171 -1745 -9115
rect -1619 -9171 -1553 -9115
rect -1427 -9171 -1361 -9115
rect -1235 -9171 -1169 -9115
rect -1043 -9171 -977 -9115
rect -851 -9171 -785 -9115
rect -659 -9171 -593 -9115
rect -467 -9171 -401 -9115
rect -275 -9171 -209 -9115
rect -83 -9171 -17 -9115
rect 109 -9171 175 -9115
rect 301 -9171 367 -9115
rect 493 -9171 559 -9115
rect 685 -9171 751 -9115
rect 877 -9171 943 -9115
rect 1069 -9171 1135 -9115
rect 1261 -9171 1327 -9115
rect 1453 -9171 1519 -9115
rect 1645 -9171 1711 -9115
rect 1837 -9171 1903 -9115
rect 2029 -9171 2095 -9115
rect 2221 -9171 2287 -9115
rect 2413 -9171 2479 -9115
rect 2605 -9171 2671 -9115
rect 2797 -9171 2863 -9115
rect 2989 -9171 3055 -9115
rect 3181 -9171 3247 -9115
rect 3373 -9171 3439 -9115
rect 3565 -9171 3631 -9115
rect 3757 -9171 3823 -9115
rect 3949 -9171 4015 -9115
rect 4141 -9171 4207 -9115
rect 4333 -9171 4399 -9115
rect 4525 -9171 4591 -9115
rect 4717 -9171 4783 -9115
rect 4909 -9171 4975 -9115
rect 5101 -9171 5167 -9115
rect 5293 -9171 5359 -9115
rect 5485 -9171 5551 -9115
rect 5691 -9181 5897 -9007
rect -4365 -10093 -4159 -9392
rect -4063 -10093 -4011 -9392
rect -4790 -11000 -4584 -10289
rect -3871 -10093 -3819 -9392
rect -3679 -10093 -3627 -9392
rect -3487 -10093 -3435 -9392
rect -3295 -10093 -3243 -9392
rect -3103 -10093 -3051 -9392
rect -2911 -10093 -2859 -9392
rect -2719 -10093 -2667 -9392
rect -2527 -10093 -2475 -9392
rect -2335 -10093 -2283 -9392
rect -2143 -10093 -2091 -9392
rect -1951 -10093 -1899 -9392
rect -1759 -10093 -1707 -9392
rect -1567 -10093 -1515 -9392
rect -1375 -10093 -1323 -9392
rect -1183 -10093 -1131 -9392
rect -991 -10093 -939 -9392
rect -799 -10093 -747 -9392
rect -607 -10093 -555 -9392
rect -415 -10093 -363 -9392
rect -223 -10093 -171 -9392
rect -31 -10093 21 -9392
rect 161 -10093 213 -9392
rect 353 -10093 405 -9392
rect 545 -10093 597 -9392
rect 737 -10093 789 -9392
rect 929 -10093 981 -9392
rect 1121 -10093 1173 -9392
rect 1313 -10093 1365 -9392
rect 1505 -10093 1557 -9392
rect 1697 -10093 1749 -9392
rect 1889 -10093 1941 -9392
rect 2081 -10093 2133 -9392
rect 2273 -10093 2325 -9392
rect 2465 -10093 2517 -9392
rect 2657 -10093 2709 -9392
rect 2849 -10093 2901 -9392
rect 3041 -10093 3093 -9392
rect 3233 -10093 3285 -9392
rect 3425 -10093 3477 -9392
rect 3617 -10093 3669 -9392
rect 3809 -10093 3861 -9392
rect 4001 -10093 4053 -9392
rect 4193 -10093 4245 -9392
rect 4385 -10093 4437 -9392
rect 4577 -10093 4629 -9392
rect 4769 -10093 4821 -9392
rect 4961 -10093 5013 -9392
rect 5153 -10093 5205 -9392
rect 5345 -10093 5397 -9392
rect 5537 -10093 5589 -9392
rect 5691 -10093 5897 -9392
rect -3971 -11000 -3905 -10289
rect -3779 -11000 -3713 -10289
rect -3587 -11000 -3521 -10289
rect -3395 -11000 -3329 -10289
rect -3203 -11000 -3137 -10289
rect -3011 -11000 -2945 -10289
rect -2819 -11000 -2753 -10289
rect -2627 -11000 -2561 -10289
rect -2435 -11000 -2369 -10289
rect -2243 -11000 -2177 -10289
rect -2051 -11000 -1985 -10289
rect -1859 -11000 -1793 -10289
rect -1667 -11000 -1601 -10289
rect -1475 -11000 -1409 -10289
rect -1283 -11000 -1217 -10289
rect -1091 -11000 -1025 -10289
rect -899 -11000 -833 -10289
rect -707 -11000 -641 -10289
rect -515 -11000 -449 -10289
rect -323 -11000 -257 -10289
rect -131 -11000 -65 -10289
rect 61 -11000 127 -10289
rect 253 -11000 319 -10289
rect 445 -11000 511 -10289
rect 637 -11000 703 -10289
rect 829 -11000 895 -10289
rect 1021 -11000 1087 -10289
rect 1213 -11000 1279 -10289
rect 1405 -11000 1471 -10289
rect 1597 -11000 1663 -10289
rect 1789 -11000 1855 -10289
rect 1981 -11000 2047 -10289
rect 2173 -11000 2239 -10289
rect 2365 -11000 2431 -10289
rect 2557 -11000 2623 -10289
rect 2749 -11000 2815 -10289
rect 2941 -11000 3007 -10289
rect 3133 -11000 3199 -10289
rect 3325 -11000 3391 -10289
rect 3517 -11000 3583 -10289
rect 3709 -11000 3775 -10289
rect 3901 -11000 3967 -10289
rect 4093 -11000 4159 -10289
rect 4285 -11000 4351 -10289
rect 4477 -11000 4543 -10289
rect 4669 -11000 4735 -10289
rect 4861 -11000 4927 -10289
rect 5053 -11000 5119 -10289
rect 5245 -11000 5311 -10289
rect 5437 -11000 5503 -10289
rect 6208 -11000 6414 -10289
rect -4365 -11399 -4159 -11225
rect -4019 -11291 -3953 -11235
rect -3827 -11291 -3761 -11235
rect -3635 -11291 -3569 -11235
rect -3443 -11291 -3377 -11235
rect -3251 -11291 -3185 -11235
rect -3059 -11291 -2993 -11235
rect -2867 -11291 -2801 -11235
rect -2675 -11291 -2609 -11235
rect -2483 -11291 -2417 -11235
rect -2291 -11291 -2225 -11235
rect -2099 -11291 -2033 -11235
rect -1907 -11291 -1841 -11235
rect -1715 -11291 -1649 -11235
rect -1523 -11291 -1457 -11235
rect -1331 -11291 -1265 -11235
rect -1139 -11291 -1073 -11235
rect -947 -11291 -881 -11235
rect -755 -11291 -689 -11235
rect -563 -11291 -497 -11235
rect -371 -11291 -305 -11235
rect -179 -11291 -113 -11235
rect 13 -11291 79 -11235
rect 205 -11291 271 -11235
rect 397 -11291 463 -11235
rect 589 -11291 655 -11235
rect 781 -11291 847 -11235
rect 973 -11291 1039 -11235
rect 1165 -11291 1231 -11235
rect 1357 -11291 1423 -11235
rect 1549 -11291 1615 -11235
rect 1741 -11291 1807 -11235
rect 1933 -11291 1999 -11235
rect 2125 -11291 2191 -11235
rect 2317 -11291 2383 -11235
rect 2509 -11291 2575 -11235
rect 2701 -11291 2767 -11235
rect 2893 -11291 2959 -11235
rect 3085 -11291 3151 -11235
rect 3277 -11291 3343 -11235
rect 3469 -11291 3535 -11235
rect 3661 -11291 3727 -11235
rect 3853 -11291 3919 -11235
rect 4045 -11291 4111 -11235
rect 4237 -11291 4303 -11235
rect 4429 -11291 4495 -11235
rect 4621 -11291 4687 -11235
rect 4813 -11291 4879 -11235
rect 5005 -11291 5071 -11235
rect 5197 -11291 5263 -11235
rect 5389 -11291 5455 -11235
rect 5691 -11399 5897 -11225
<< metal2 >>
rect 29 1715 1503 2262
rect 2398 1715 4108 1725
rect -2576 1435 383 1715
rect 441 1435 855 1715
rect 913 1435 1327 1715
rect 1385 1435 2408 1715
rect -2576 1415 -144 1435
rect 383 1425 441 1435
rect 855 1425 913 1435
rect 1327 1425 1385 1435
rect 1676 1425 2408 1435
rect 4098 1425 4108 1715
rect 1676 1415 4108 1425
rect -4849 1369 6391 1379
rect -4849 1076 -3193 1369
rect -2900 1366 4442 1369
rect -2900 1076 29 1366
rect -4849 1066 29 1076
rect 87 1066 265 1366
rect 323 1066 501 1366
rect 559 1066 737 1366
rect 795 1066 973 1366
rect 1031 1066 1209 1366
rect 1267 1066 1445 1366
rect 1503 1076 4442 1366
rect 4735 1076 6391 1369
rect 1503 1066 6391 1076
rect 29 1056 87 1066
rect 265 1056 323 1066
rect 501 1056 559 1066
rect 737 1056 795 1066
rect 973 1056 1031 1066
rect 1209 1056 1267 1066
rect 1445 1056 1503 1066
rect 147 1015 205 1025
rect 619 1015 677 1025
rect 1091 1015 1149 1025
rect -2576 1005 147 1015
rect -2576 725 -2566 1005
rect -876 725 147 1005
rect -2576 715 147 725
rect 205 715 619 1015
rect 677 715 1091 1015
rect 1149 715 4108 1015
rect 147 705 205 715
rect 619 705 677 715
rect 1091 705 1149 715
rect -4849 225 6472 387
rect -4849 69 321 225
rect 1211 69 6472 225
rect 321 59 1211 69
rect -2678 -202 -2619 -192
rect -823 -202 -764 -192
rect -2619 -268 -823 -202
rect -2678 -278 -2619 -268
rect -823 -278 -764 -268
rect -2576 -309 -2222 -299
rect -2164 -309 -1750 -299
rect -1692 -309 -1278 -299
rect -1220 -309 -866 -299
rect -2576 -589 -2566 -309
rect -876 -589 -866 -309
rect -2576 -599 -2222 -589
rect -2164 -599 -1750 -589
rect -1692 -599 -1278 -589
rect -1220 -599 -866 -589
rect -2222 -609 -2164 -599
rect -1750 -609 -1692 -599
rect -1278 -609 -1220 -599
rect -2678 -649 -2619 -639
rect -2458 -649 -2400 -639
rect -1986 -649 -1928 -639
rect -1514 -649 -1456 -639
rect -1042 -649 -984 -639
rect -823 -649 -764 -639
rect -617 -649 -317 8
rect -63 -18 2149 8
rect -63 -472 421 -18
rect 479 -472 1053 -18
rect 1111 -472 2149 -18
rect 2296 -202 2355 -192
rect 4151 -202 4210 -192
rect 2355 -268 4151 -202
rect 2296 -278 2355 -268
rect 4151 -278 4210 -268
rect -2619 -949 -2458 -649
rect -2400 -949 -1986 -649
rect -1928 -949 -1514 -649
rect -1456 -949 -1042 -649
rect -984 -949 -823 -649
rect -764 -949 -317 -649
rect -2678 -959 -2619 -949
rect -2458 -959 -2400 -949
rect -1986 -959 -1928 -949
rect -1514 -959 -1456 -949
rect -1042 -959 -984 -949
rect -823 -959 -764 -949
rect -2576 -999 -2518 -989
rect -2340 -999 -2282 -989
rect -2104 -999 -2046 -989
rect -1868 -999 -1810 -989
rect -1632 -999 -1574 -989
rect -1396 -999 -1338 -989
rect -1160 -999 -1102 -989
rect -924 -999 -866 -989
rect -2668 -1009 -2576 -999
rect -2518 -1009 -2340 -999
rect -2282 -1009 -2104 -999
rect -2046 -1009 -1868 -999
rect -1810 -1009 -1632 -999
rect -1574 -1009 -1396 -999
rect -1338 -1009 -1160 -999
rect -1102 -1009 -924 -999
rect -2668 -1299 -2576 -1289
rect -2518 -1299 -2340 -1289
rect -2282 -1299 -2104 -1289
rect -2046 -1299 -1868 -1289
rect -1810 -1299 -1632 -1289
rect -1574 -1299 -1396 -1289
rect -1338 -1299 -1160 -1289
rect -1102 -1299 -924 -1289
rect -2576 -1309 -2518 -1299
rect -924 -1309 -866 -1299
rect -617 -1145 -317 -949
rect -63 -1090 -53 -527
rect 5 -537 263 -527
rect 321 -537 579 -527
rect 394 -1080 579 -537
rect 5 -1090 263 -1080
rect 321 -1090 579 -1080
rect 637 -1090 895 -527
rect 953 -537 1211 -527
rect 1269 -537 1527 -527
rect 953 -1080 1138 -537
rect 953 -1090 1211 -1080
rect 1269 -1090 1527 -1080
rect 1585 -1090 1595 -527
rect 1849 -649 2149 -472
rect 2398 -309 2752 -299
rect 2810 -309 3224 -299
rect 3282 -309 3696 -299
rect 3754 -309 4108 -299
rect 2398 -589 2408 -309
rect 4098 -589 4108 -309
rect 2398 -599 2752 -589
rect 2810 -599 3224 -589
rect 3282 -599 3696 -589
rect 3754 -599 4108 -589
rect 2752 -609 2810 -599
rect 3224 -609 3282 -599
rect 3696 -609 3754 -599
rect 2296 -649 2355 -639
rect 2516 -649 2574 -639
rect 2988 -649 3046 -639
rect 3460 -649 3518 -639
rect 3932 -649 3990 -639
rect 4151 -649 4210 -639
rect 1849 -949 2296 -649
rect 2355 -949 2516 -649
rect 2574 -949 2988 -649
rect 3046 -949 3460 -649
rect 3518 -949 3932 -649
rect 3990 -949 4151 -649
rect 737 -1145 795 -1135
rect -2678 -1337 -2619 -1327
rect -2403 -1337 -1039 -1327
rect -823 -1337 -764 -1327
rect -2619 -1396 -2403 -1337
rect -1039 -1396 -823 -1337
rect -2678 -1406 -2619 -1396
rect -2403 -1406 -1039 -1396
rect -823 -1406 -764 -1396
rect -617 -1599 105 -1145
rect 163 -1599 737 -1145
rect 795 -1599 1369 -1145
rect 1427 -1599 1595 -1145
rect -617 -1625 1595 -1599
rect 1849 -1625 2149 -949
rect 2296 -959 2355 -949
rect 2516 -959 2574 -949
rect 2988 -959 3046 -949
rect 3460 -959 3518 -949
rect 3932 -959 3990 -949
rect 4151 -959 4210 -949
rect 2398 -999 2456 -989
rect 2634 -999 2692 -989
rect 2870 -999 2928 -989
rect 3106 -999 3164 -989
rect 3342 -999 3400 -989
rect 3578 -999 3636 -989
rect 3814 -999 3872 -989
rect 4050 -999 4108 -989
rect 2456 -1009 2634 -999
rect 2692 -1009 2870 -999
rect 2928 -1009 3106 -999
rect 3164 -1009 3342 -999
rect 3400 -1009 3578 -999
rect 3636 -1009 3814 -999
rect 3872 -1009 4050 -999
rect 4108 -1009 4201 -999
rect 2456 -1299 2634 -1289
rect 2692 -1299 2870 -1289
rect 2928 -1299 3106 -1289
rect 3164 -1299 3342 -1289
rect 3400 -1299 3578 -1289
rect 3636 -1299 3814 -1289
rect 3872 -1299 4050 -1289
rect 4108 -1299 4201 -1289
rect 2398 -1309 2456 -1299
rect 4050 -1309 4108 -1299
rect 2296 -1337 2355 -1327
rect 2571 -1337 3935 -1327
rect 4151 -1337 4210 -1327
rect 2355 -1396 2571 -1337
rect 3935 -1396 4151 -1337
rect 2296 -1406 2355 -1396
rect 2571 -1406 3935 -1396
rect 4151 -1406 4210 -1396
rect 163 -1667 1369 -1657
rect -4849 -1823 163 -1667
rect 1369 -1823 6472 -1667
rect -4849 -1985 6472 -1823
rect -1942 -2382 3484 -2372
rect -1942 -2597 -1932 -2382
rect -1707 -2597 -1259 -2382
rect -1942 -2607 -1259 -2597
rect 2791 -2388 3484 -2382
rect 2791 -2603 3249 -2388
rect 3474 -2603 3484 -2388
rect 2791 -2607 3484 -2603
rect -1269 -2617 3484 -2607
rect -1585 -2655 3117 -2645
rect -1585 -2948 -1327 -2655
rect -1269 -2948 -1132 -2655
rect -688 -2948 -295 -2655
rect -237 -2948 -50 -2655
rect 394 -2948 737 -2655
rect 795 -2948 1138 -2655
rect 1582 -2948 1769 -2655
rect 1827 -2948 2220 -2655
rect 2664 -2948 2801 -2655
rect 2859 -2948 3117 -2655
rect -1585 -2958 3117 -2948
rect -4781 -2996 6472 -2986
rect -4781 -3294 -1932 -2996
rect -1707 -3294 -811 -2996
rect -753 -3294 221 -2996
rect 279 -3294 1253 -2996
rect 1311 -3294 2285 -2996
rect 2343 -3294 3249 -2996
rect 3474 -3294 6472 -2996
rect -4781 -3304 6472 -3294
rect -3203 -3342 -2091 -3332
rect -3203 -3635 -3193 -3342
rect -2900 -3635 -2091 -3342
rect -3203 -3645 -2091 -3635
rect -2001 -3342 3543 -3332
rect -2001 -3635 -1585 -3342
rect -1527 -3635 -1069 -3342
rect -1011 -3635 -593 -3342
rect -149 -3635 -37 -3342
rect 21 -3635 479 -3342
rect 537 -3635 995 -3342
rect 1053 -3635 1511 -3342
rect 1569 -3635 1677 -3342
rect 2121 -3635 2543 -3342
rect 2601 -3635 3059 -3342
rect 3117 -3635 3543 -3342
rect -2001 -3645 3543 -3635
rect 3633 -3342 4745 -3332
rect 3633 -3635 4442 -3342
rect 4735 -3635 4745 -3342
rect 3633 -3645 4745 -3635
rect -1932 -3683 3249 -3673
rect -1707 -3908 -1259 -3683
rect 2791 -3693 3474 -3683
rect 2791 -3908 3249 -3693
rect -1932 -3918 3474 -3908
rect -4791 -4262 -4584 -4252
rect 6208 -4262 6415 -4252
rect -4584 -4272 6208 -4262
rect -4584 -4425 -1132 -4272
rect -688 -4425 -50 -4272
rect 394 -4425 1138 -4272
rect 1582 -4425 2220 -4272
rect 2664 -4425 6208 -4272
rect -4584 -4435 6208 -4425
rect -4791 -4445 -4584 -4435
rect 6208 -4445 6415 -4435
rect -4974 -4571 -4841 -4561
rect -4365 -4571 -4159 -4561
rect 5691 -4571 5897 -4561
rect 6465 -4571 6598 -4561
rect -4841 -4745 -4365 -4571
rect -4159 -4581 5691 -4571
rect -4159 -4679 -593 -4581
rect -149 -4679 1677 -4581
rect 2121 -4679 5691 -4581
rect -4159 -4735 -3923 -4679
rect -3857 -4735 -3731 -4679
rect -3665 -4735 -3539 -4679
rect -3473 -4735 -3347 -4679
rect -3281 -4735 -3155 -4679
rect -3089 -4735 -2963 -4679
rect -2897 -4735 -2771 -4679
rect -2705 -4735 -2579 -4679
rect -2513 -4735 -2387 -4679
rect -2321 -4735 -2195 -4679
rect -2129 -4735 -2003 -4679
rect -1937 -4735 -1811 -4679
rect -1745 -4735 -1619 -4679
rect -1553 -4735 -1427 -4679
rect -1361 -4735 -1235 -4679
rect -1169 -4735 -1043 -4679
rect -977 -4735 -851 -4679
rect -785 -4735 -659 -4679
rect -149 -4735 -83 -4679
rect -17 -4735 109 -4679
rect 175 -4735 301 -4679
rect 367 -4735 493 -4679
rect 559 -4735 685 -4679
rect 751 -4735 877 -4679
rect 943 -4735 1069 -4679
rect 1135 -4735 1261 -4679
rect 1327 -4735 1453 -4679
rect 1519 -4735 1645 -4679
rect 2121 -4735 2221 -4679
rect 2287 -4735 2413 -4679
rect 2479 -4735 2605 -4679
rect 2671 -4735 2797 -4679
rect 2863 -4735 2989 -4679
rect 3055 -4735 3181 -4679
rect 3247 -4735 3373 -4679
rect 3439 -4735 3565 -4679
rect 3631 -4735 3757 -4679
rect 3823 -4735 3949 -4679
rect 4015 -4735 4141 -4679
rect 4207 -4735 4333 -4679
rect 4399 -4735 4525 -4679
rect 4591 -4735 4717 -4679
rect 4783 -4735 4909 -4679
rect 4975 -4735 5101 -4679
rect 5167 -4735 5293 -4679
rect 5359 -4735 5485 -4679
rect 5551 -4735 5691 -4679
rect -4159 -4745 5691 -4735
rect 5897 -4745 6465 -4571
rect -4841 -4956 6465 -4745
rect -4841 -5657 -4365 -4956
rect -4159 -5657 -4063 -4956
rect -4011 -5657 -3871 -4956
rect -3819 -5657 -3679 -4956
rect -3627 -5657 -3487 -4956
rect -3435 -5657 -3295 -4956
rect -3243 -5657 -3103 -4956
rect -3051 -5657 -2911 -4956
rect -2859 -5657 -2719 -4956
rect -2667 -5657 -2527 -4956
rect -2475 -5657 -2335 -4956
rect -2283 -5657 -2143 -4956
rect -2091 -5657 -1951 -4956
rect -1899 -5657 -1759 -4956
rect -1707 -5657 -1567 -4956
rect -1515 -5657 -1375 -4956
rect -1323 -5657 -1183 -4956
rect -1131 -5657 -991 -4956
rect -939 -5657 -799 -4956
rect -747 -5657 -607 -4956
rect -555 -5657 -415 -4956
rect -363 -5657 -223 -4956
rect -171 -5657 -31 -4956
rect 21 -5657 161 -4956
rect 213 -5657 353 -4956
rect 405 -5657 545 -4956
rect 597 -5657 737 -4956
rect 789 -5657 929 -4956
rect 981 -5657 1121 -4956
rect 1173 -5657 1313 -4956
rect 1365 -5657 1505 -4956
rect 1557 -5657 1697 -4956
rect 1749 -5657 1889 -4956
rect 1941 -5657 2081 -4956
rect 2133 -5657 2273 -4956
rect 2325 -5657 2465 -4956
rect 2517 -5657 2657 -4956
rect 2709 -5657 2849 -4956
rect 2901 -5657 3041 -4956
rect 3093 -5657 3233 -4956
rect 3285 -5657 3425 -4956
rect 3477 -5657 3617 -4956
rect 3669 -5657 3809 -4956
rect 3861 -5657 4001 -4956
rect 4053 -5657 4193 -4956
rect 4245 -5657 4385 -4956
rect 4437 -5657 4577 -4956
rect 4629 -5657 4769 -4956
rect 4821 -5657 4961 -4956
rect 5013 -5657 5153 -4956
rect 5205 -5657 5345 -4956
rect 5397 -5657 5537 -4956
rect 5589 -5657 5691 -4956
rect 5897 -5657 6465 -4956
rect -4974 -5667 -4841 -5657
rect -4365 -5667 -4159 -5657
rect 5537 -5667 5589 -5657
rect 5691 -5667 5897 -5657
rect 6465 -5667 6598 -5657
rect -4790 -5853 -4584 -5843
rect 6208 -5853 6414 -5843
rect -4584 -6564 -3971 -5853
rect -3905 -6564 -3779 -5853
rect -3713 -6564 -3587 -5853
rect -3521 -6564 -3395 -5853
rect -3329 -6564 -3203 -5853
rect -3137 -6564 -3011 -5853
rect -2945 -6564 -2819 -5853
rect -2753 -6564 -2627 -5853
rect -2561 -6564 -2435 -5853
rect -2369 -6564 -2243 -5853
rect -2177 -6564 -2051 -5853
rect -1985 -6564 -1859 -5853
rect -1793 -6564 -1667 -5853
rect -1601 -6564 -1475 -5853
rect -1409 -6564 -1283 -5853
rect -1217 -6564 -1091 -5853
rect -1025 -6564 -899 -5853
rect -833 -6564 -707 -5853
rect -641 -6564 -515 -5853
rect -449 -6564 -323 -5853
rect -257 -6564 -131 -5853
rect -65 -6564 61 -5853
rect 127 -6564 253 -5853
rect 319 -6564 445 -5853
rect 511 -6564 637 -5853
rect 703 -6564 829 -5853
rect 895 -6564 1021 -5853
rect 1087 -6564 1213 -5853
rect 1279 -6564 1405 -5853
rect 1471 -6564 1597 -5853
rect 1663 -6564 1789 -5853
rect 1855 -6564 1981 -5853
rect 2047 -6564 2173 -5853
rect 2239 -6564 2365 -5853
rect 2431 -6564 2557 -5853
rect 2623 -6564 2749 -5853
rect 2815 -6564 2941 -5853
rect 3007 -6564 3133 -5853
rect 3199 -6564 3325 -5853
rect 3391 -6564 3517 -5853
rect 3583 -6564 3709 -5853
rect 3775 -6564 3901 -5853
rect 3967 -6564 4093 -5853
rect 4159 -6564 4285 -5853
rect 4351 -6564 4477 -5853
rect 4543 -6564 4669 -5853
rect 4735 -6564 4861 -5853
rect 4927 -6564 5053 -5853
rect 5119 -6564 5245 -5853
rect 5311 -6564 5437 -5853
rect 5503 -6564 6208 -5853
rect -4790 -6574 -4584 -6564
rect 6208 -6574 6414 -6564
rect -4365 -6789 -4159 -6779
rect 5691 -6789 5897 -6779
rect -4159 -6799 5691 -6789
rect -4159 -6855 -4019 -6799
rect -3953 -6855 -3827 -6799
rect -3761 -6855 -3635 -6799
rect -3569 -6855 -3443 -6799
rect -3377 -6855 -3251 -6799
rect -3185 -6855 -3059 -6799
rect -2993 -6855 -2867 -6799
rect -2801 -6855 -2675 -6799
rect -2609 -6855 -2483 -6799
rect -2417 -6855 -2291 -6799
rect -2225 -6855 -2099 -6799
rect -2033 -6855 -1907 -6799
rect -1841 -6855 -1715 -6799
rect -1649 -6855 -1523 -6799
rect -1457 -6855 -1331 -6799
rect -1265 -6855 -1139 -6799
rect -1073 -6855 -947 -6799
rect -881 -6855 -755 -6799
rect -689 -6855 -563 -6799
rect -497 -6855 -371 -6799
rect -305 -6855 -179 -6799
rect -113 -6855 13 -6799
rect 79 -6855 205 -6799
rect 271 -6855 397 -6799
rect 463 -6855 589 -6799
rect 655 -6855 781 -6799
rect 847 -6855 973 -6799
rect 1039 -6855 1165 -6799
rect 1231 -6855 1357 -6799
rect 1423 -6855 1549 -6799
rect 1615 -6855 1741 -6799
rect 1807 -6855 1933 -6799
rect 1999 -6855 2125 -6799
rect 2191 -6855 2317 -6799
rect 2383 -6855 2509 -6799
rect 2575 -6855 2701 -6799
rect 2767 -6855 2893 -6799
rect 2959 -6855 3085 -6799
rect 3151 -6855 3277 -6799
rect 3343 -6855 3469 -6799
rect 3535 -6855 3661 -6799
rect 3727 -6855 3853 -6799
rect 3919 -6855 4045 -6799
rect 4111 -6855 4237 -6799
rect 4303 -6855 4429 -6799
rect 4495 -6855 4621 -6799
rect 4687 -6855 4813 -6799
rect 4879 -6855 5005 -6799
rect 5071 -6855 5197 -6799
rect 5263 -6855 5389 -6799
rect 5455 -6855 5691 -6799
rect -4159 -6897 5691 -6855
rect -4159 -6953 -4019 -6897
rect -3953 -6953 -3827 -6897
rect -3761 -6953 -3635 -6897
rect -3569 -6953 -3443 -6897
rect -3377 -6953 -3251 -6897
rect -3185 -6953 -3059 -6897
rect -2993 -6953 -2867 -6897
rect -2801 -6953 -2675 -6897
rect -2609 -6953 -2483 -6897
rect -2417 -6953 -2291 -6897
rect -2225 -6953 -2099 -6897
rect -2033 -6953 -1907 -6897
rect -1841 -6953 -1715 -6897
rect -1649 -6953 -1523 -6897
rect -1457 -6953 -1331 -6897
rect -1265 -6953 -1139 -6897
rect -1073 -6953 -947 -6897
rect -881 -6953 -755 -6897
rect -689 -6953 -563 -6897
rect -497 -6953 -371 -6897
rect -305 -6953 -179 -6897
rect -113 -6953 13 -6897
rect 79 -6953 205 -6897
rect 271 -6953 397 -6897
rect 463 -6953 589 -6897
rect 655 -6953 781 -6897
rect 847 -6953 973 -6897
rect 1039 -6953 1165 -6897
rect 1231 -6953 1357 -6897
rect 1423 -6953 1549 -6897
rect 1615 -6953 1741 -6897
rect 1807 -6953 1933 -6897
rect 1999 -6953 2125 -6897
rect 2191 -6953 2317 -6897
rect 2383 -6953 2509 -6897
rect 2575 -6953 2701 -6897
rect 2767 -6953 2893 -6897
rect 2959 -6953 3085 -6897
rect 3151 -6953 3277 -6897
rect 3343 -6953 3469 -6897
rect 3535 -6953 3661 -6897
rect 3727 -6953 3853 -6897
rect 3919 -6953 4045 -6897
rect 4111 -6953 4237 -6897
rect 4303 -6953 4429 -6897
rect 4495 -6953 4621 -6897
rect 4687 -6953 4813 -6897
rect 4879 -6953 5005 -6897
rect 5071 -6953 5197 -6897
rect 5263 -6953 5389 -6897
rect 5455 -6953 5691 -6897
rect -4159 -6963 5691 -6953
rect -4365 -6973 -4159 -6963
rect 5691 -6973 5897 -6963
rect -4365 -7174 -4159 -7164
rect 5537 -7174 5589 -7164
rect 5691 -7174 5897 -7164
rect -4159 -7875 -4063 -7174
rect -4011 -7875 -3871 -7174
rect -3819 -7875 -3679 -7174
rect -3627 -7875 -3487 -7174
rect -3435 -7875 -3295 -7174
rect -3243 -7875 -3103 -7174
rect -3051 -7875 -2911 -7174
rect -2859 -7875 -2719 -7174
rect -2667 -7875 -2527 -7174
rect -2475 -7875 -2335 -7174
rect -2283 -7875 -2143 -7174
rect -2091 -7875 -1951 -7174
rect -1899 -7875 -1759 -7174
rect -1707 -7875 -1567 -7174
rect -1515 -7875 -1375 -7174
rect -1323 -7875 -1183 -7174
rect -1131 -7875 -991 -7174
rect -939 -7875 -799 -7174
rect -747 -7875 -607 -7174
rect -555 -7875 -415 -7174
rect -363 -7875 -223 -7174
rect -171 -7875 -31 -7174
rect 21 -7875 161 -7174
rect 213 -7875 353 -7174
rect 405 -7875 545 -7174
rect 597 -7875 737 -7174
rect 789 -7875 929 -7174
rect 981 -7875 1121 -7174
rect 1173 -7875 1313 -7174
rect 1365 -7875 1505 -7174
rect 1557 -7875 1697 -7174
rect 1749 -7875 1889 -7174
rect 1941 -7875 2081 -7174
rect 2133 -7875 2273 -7174
rect 2325 -7875 2465 -7174
rect 2517 -7875 2657 -7174
rect 2709 -7875 2849 -7174
rect 2901 -7875 3041 -7174
rect 3093 -7875 3233 -7174
rect 3285 -7875 3425 -7174
rect 3477 -7875 3617 -7174
rect 3669 -7875 3809 -7174
rect 3861 -7875 4001 -7174
rect 4053 -7875 4193 -7174
rect 4245 -7875 4385 -7174
rect 4437 -7875 4577 -7174
rect 4629 -7875 4769 -7174
rect 4821 -7875 4961 -7174
rect 5013 -7875 5153 -7174
rect 5205 -7875 5345 -7174
rect 5397 -7875 5537 -7174
rect 5589 -7875 5691 -7174
rect -4365 -7885 -4159 -7875
rect 5537 -7885 5589 -7875
rect 5691 -7885 5897 -7875
rect -4790 -8071 -4584 -8061
rect 6208 -8071 6414 -8061
rect -4584 -8782 -3971 -8071
rect -3905 -8782 -3779 -8071
rect -3713 -8782 -3587 -8071
rect -3521 -8782 -3395 -8071
rect -3329 -8782 -3203 -8071
rect -3137 -8782 -3011 -8071
rect -2945 -8782 -2819 -8071
rect -2753 -8782 -2627 -8071
rect -2561 -8782 -2435 -8071
rect -2369 -8782 -2243 -8071
rect -2177 -8782 -2051 -8071
rect -1985 -8782 -1859 -8071
rect -1793 -8782 -1667 -8071
rect -1601 -8782 -1475 -8071
rect -1409 -8782 -1283 -8071
rect -1217 -8782 -1091 -8071
rect -1025 -8782 -899 -8071
rect -833 -8782 -707 -8071
rect -641 -8782 -515 -8071
rect -449 -8782 -323 -8071
rect -257 -8782 -131 -8071
rect -65 -8782 61 -8071
rect 127 -8782 253 -8071
rect 319 -8782 445 -8071
rect 511 -8782 637 -8071
rect 703 -8782 829 -8071
rect 895 -8782 1021 -8071
rect 1087 -8782 1213 -8071
rect 1279 -8782 1405 -8071
rect 1471 -8782 1597 -8071
rect 1663 -8782 1789 -8071
rect 1855 -8782 1981 -8071
rect 2047 -8782 2173 -8071
rect 2239 -8782 2365 -8071
rect 2431 -8782 2557 -8071
rect 2623 -8782 2749 -8071
rect 2815 -8782 2941 -8071
rect 3007 -8782 3133 -8071
rect 3199 -8782 3325 -8071
rect 3391 -8782 3517 -8071
rect 3583 -8782 3709 -8071
rect 3775 -8782 3901 -8071
rect 3967 -8782 4093 -8071
rect 4159 -8782 4285 -8071
rect 4351 -8782 4477 -8071
rect 4543 -8782 4669 -8071
rect 4735 -8782 4861 -8071
rect 4927 -8782 5053 -8071
rect 5119 -8782 5245 -8071
rect 5311 -8782 5437 -8071
rect 5503 -8782 6208 -8071
rect -4790 -8792 -4584 -8782
rect 6208 -8792 6414 -8782
rect -4365 -9007 -4159 -8997
rect 5691 -9007 5897 -8997
rect -4365 -9017 5691 -9007
rect -4365 -9071 -3923 -9017
rect -4159 -9073 -3923 -9071
rect -3857 -9073 -3731 -9017
rect -3665 -9073 -3539 -9017
rect -3473 -9073 -3347 -9017
rect -3281 -9073 -3155 -9017
rect -3089 -9073 -2963 -9017
rect -2897 -9073 -2771 -9017
rect -2705 -9073 -2579 -9017
rect -2513 -9073 -2387 -9017
rect -2321 -9073 -2195 -9017
rect -2129 -9073 -2003 -9017
rect -1937 -9073 -1811 -9017
rect -1745 -9073 -1619 -9017
rect -1553 -9073 -1427 -9017
rect -1361 -9073 -1235 -9017
rect -1169 -9073 -1043 -9017
rect -977 -9073 -851 -9017
rect -785 -9073 -659 -9017
rect -593 -9073 -467 -9017
rect -401 -9073 -275 -9017
rect -209 -9073 -83 -9017
rect -17 -9073 109 -9017
rect 175 -9073 301 -9017
rect 367 -9073 493 -9017
rect 559 -9073 685 -9017
rect 751 -9073 877 -9017
rect 943 -9073 1069 -9017
rect 1135 -9073 1261 -9017
rect 1327 -9073 1453 -9017
rect 1519 -9073 1645 -9017
rect 1711 -9073 1837 -9017
rect 1903 -9073 2029 -9017
rect 2095 -9073 2221 -9017
rect 2287 -9073 2413 -9017
rect 2479 -9073 2605 -9017
rect 2671 -9073 2797 -9017
rect 2863 -9073 2989 -9017
rect 3055 -9073 3181 -9017
rect 3247 -9073 3373 -9017
rect 3439 -9073 3565 -9017
rect 3631 -9073 3757 -9017
rect 3823 -9073 3949 -9017
rect 4015 -9073 4141 -9017
rect 4207 -9073 4333 -9017
rect 4399 -9073 4525 -9017
rect 4591 -9073 4717 -9017
rect 4783 -9073 4909 -9017
rect 4975 -9073 5101 -9017
rect 5167 -9073 5293 -9017
rect 5359 -9073 5485 -9017
rect 5551 -9073 5691 -9017
rect -4159 -9115 5691 -9073
rect -4159 -9171 -3923 -9115
rect -3857 -9171 -3731 -9115
rect -3665 -9171 -3539 -9115
rect -3473 -9171 -3347 -9115
rect -3281 -9171 -3155 -9115
rect -3089 -9171 -2963 -9115
rect -2897 -9171 -2771 -9115
rect -2705 -9171 -2579 -9115
rect -2513 -9171 -2387 -9115
rect -2321 -9171 -2195 -9115
rect -2129 -9171 -2003 -9115
rect -1937 -9171 -1811 -9115
rect -1745 -9171 -1619 -9115
rect -1553 -9171 -1427 -9115
rect -1361 -9171 -1235 -9115
rect -1169 -9171 -1043 -9115
rect -977 -9171 -851 -9115
rect -785 -9171 -659 -9115
rect -593 -9171 -467 -9115
rect -401 -9171 -275 -9115
rect -209 -9171 -83 -9115
rect -17 -9171 109 -9115
rect 175 -9171 301 -9115
rect 367 -9171 493 -9115
rect 559 -9171 685 -9115
rect 751 -9171 877 -9115
rect 943 -9171 1069 -9115
rect 1135 -9171 1261 -9115
rect 1327 -9171 1453 -9115
rect 1519 -9171 1645 -9115
rect 1711 -9171 1837 -9115
rect 1903 -9171 2029 -9115
rect 2095 -9171 2221 -9115
rect 2287 -9171 2413 -9115
rect 2479 -9171 2605 -9115
rect 2671 -9171 2797 -9115
rect 2863 -9171 2989 -9115
rect 3055 -9171 3181 -9115
rect 3247 -9171 3373 -9115
rect 3439 -9171 3565 -9115
rect 3631 -9171 3757 -9115
rect 3823 -9171 3949 -9115
rect 4015 -9171 4141 -9115
rect 4207 -9171 4333 -9115
rect 4399 -9171 4525 -9115
rect 4591 -9171 4717 -9115
rect 4783 -9171 4909 -9115
rect 4975 -9171 5101 -9115
rect 5167 -9171 5293 -9115
rect 5359 -9171 5485 -9115
rect 5551 -9171 5691 -9115
rect -4159 -9181 5691 -9171
rect -4365 -9191 -4159 -9181
rect 5691 -9191 5897 -9181
rect -4365 -9392 -4159 -9382
rect 5537 -9392 5589 -9382
rect 5691 -9392 5897 -9382
rect -4159 -10093 -4063 -9392
rect -4011 -10093 -3871 -9392
rect -3819 -10093 -3679 -9392
rect -3627 -10093 -3487 -9392
rect -3435 -10093 -3295 -9392
rect -3243 -10093 -3103 -9392
rect -3051 -10093 -2911 -9392
rect -2859 -10093 -2719 -9392
rect -2667 -10093 -2527 -9392
rect -2475 -10093 -2335 -9392
rect -2283 -10093 -2143 -9392
rect -2091 -10093 -1951 -9392
rect -1899 -10093 -1759 -9392
rect -1707 -10093 -1567 -9392
rect -1515 -10093 -1375 -9392
rect -1323 -10093 -1183 -9392
rect -1131 -10093 -991 -9392
rect -939 -10093 -799 -9392
rect -747 -10093 -607 -9392
rect -555 -10093 -415 -9392
rect -363 -10093 -223 -9392
rect -171 -10093 -31 -9392
rect 21 -10093 161 -9392
rect 213 -10093 353 -9392
rect 405 -10093 545 -9392
rect 597 -10093 737 -9392
rect 789 -10093 929 -9392
rect 981 -10093 1121 -9392
rect 1173 -10093 1313 -9392
rect 1365 -10093 1505 -9392
rect 1557 -10093 1697 -9392
rect 1749 -10093 1889 -9392
rect 1941 -10093 2081 -9392
rect 2133 -10093 2273 -9392
rect 2325 -10093 2465 -9392
rect 2517 -10093 2657 -9392
rect 2709 -10093 2849 -9392
rect 2901 -10093 3041 -9392
rect 3093 -10093 3233 -9392
rect 3285 -10093 3425 -9392
rect 3477 -10093 3617 -9392
rect 3669 -10093 3809 -9392
rect 3861 -10093 4001 -9392
rect 4053 -10093 4193 -9392
rect 4245 -10093 4385 -9392
rect 4437 -10093 4577 -9392
rect 4629 -10093 4769 -9392
rect 4821 -10093 4961 -9392
rect 5013 -10093 5153 -9392
rect 5205 -10093 5345 -9392
rect 5397 -10093 5537 -9392
rect 5589 -10093 5691 -9392
rect -4365 -10103 -4159 -10093
rect 5537 -10103 5589 -10093
rect 5691 -10103 5897 -10093
rect -4790 -10289 -4584 -10279
rect 6208 -10289 6414 -10279
rect -4584 -11000 -3971 -10289
rect -3905 -11000 -3779 -10289
rect -3713 -11000 -3587 -10289
rect -3521 -11000 -3395 -10289
rect -3329 -11000 -3203 -10289
rect -3137 -11000 -3011 -10289
rect -2945 -11000 -2819 -10289
rect -2753 -11000 -2627 -10289
rect -2561 -11000 -2435 -10289
rect -2369 -11000 -2243 -10289
rect -2177 -11000 -2051 -10289
rect -1985 -11000 -1859 -10289
rect -1793 -11000 -1667 -10289
rect -1601 -11000 -1475 -10289
rect -1409 -11000 -1283 -10289
rect -1217 -11000 -1091 -10289
rect -1025 -11000 -899 -10289
rect -833 -11000 -707 -10289
rect -641 -11000 -515 -10289
rect -449 -11000 -323 -10289
rect -257 -11000 -131 -10289
rect -65 -11000 61 -10289
rect 127 -11000 253 -10289
rect 319 -11000 445 -10289
rect 511 -11000 637 -10289
rect 703 -11000 829 -10289
rect 895 -11000 1021 -10289
rect 1087 -11000 1213 -10289
rect 1279 -11000 1405 -10289
rect 1471 -11000 1597 -10289
rect 1663 -11000 1789 -10289
rect 1855 -11000 1981 -10289
rect 2047 -11000 2173 -10289
rect 2239 -11000 2365 -10289
rect 2431 -11000 2557 -10289
rect 2623 -11000 2749 -10289
rect 2815 -11000 2941 -10289
rect 3007 -11000 3133 -10289
rect 3199 -11000 3325 -10289
rect 3391 -11000 3517 -10289
rect 3583 -11000 3709 -10289
rect 3775 -11000 3901 -10289
rect 3967 -11000 4093 -10289
rect 4159 -11000 4285 -10289
rect 4351 -11000 4477 -10289
rect 4543 -11000 4669 -10289
rect 4735 -11000 4861 -10289
rect 4927 -11000 5053 -10289
rect 5119 -11000 5245 -10289
rect 5311 -11000 5437 -10289
rect 5503 -11000 6208 -10289
rect -4790 -11010 -4584 -11000
rect 6208 -11010 6414 -11000
rect -4365 -11225 -4159 -11215
rect 5691 -11225 5897 -11215
rect -4159 -11235 5691 -11225
rect -4159 -11291 -4019 -11235
rect -3953 -11291 -3827 -11235
rect -3761 -11291 -3635 -11235
rect -3569 -11291 -3443 -11235
rect -3377 -11291 -3251 -11235
rect -3185 -11291 -3059 -11235
rect -2993 -11291 -2867 -11235
rect -2801 -11291 -2675 -11235
rect -2609 -11291 -2483 -11235
rect -2417 -11291 -2291 -11235
rect -2225 -11291 -2099 -11235
rect -2033 -11291 -1907 -11235
rect -1841 -11291 -1715 -11235
rect -1649 -11291 -1523 -11235
rect -1457 -11291 -1331 -11235
rect -1265 -11291 -1139 -11235
rect -1073 -11291 -947 -11235
rect -881 -11291 -755 -11235
rect -689 -11291 -563 -11235
rect -497 -11291 -371 -11235
rect -305 -11291 -179 -11235
rect -113 -11291 13 -11235
rect 79 -11291 205 -11235
rect 271 -11291 397 -11235
rect 463 -11291 589 -11235
rect 655 -11291 781 -11235
rect 847 -11291 973 -11235
rect 1039 -11291 1165 -11235
rect 1231 -11291 1357 -11235
rect 1423 -11291 1549 -11235
rect 1615 -11291 1741 -11235
rect 1807 -11291 1933 -11235
rect 1999 -11291 2125 -11235
rect 2191 -11291 2317 -11235
rect 2383 -11291 2509 -11235
rect 2575 -11291 2701 -11235
rect 2767 -11291 2893 -11235
rect 2959 -11291 3085 -11235
rect 3151 -11291 3277 -11235
rect 3343 -11291 3469 -11235
rect 3535 -11291 3661 -11235
rect 3727 -11291 3853 -11235
rect 3919 -11291 4045 -11235
rect 4111 -11291 4237 -11235
rect 4303 -11291 4429 -11235
rect 4495 -11291 4621 -11235
rect 4687 -11291 4813 -11235
rect 4879 -11291 5005 -11235
rect 5071 -11291 5197 -11235
rect 5263 -11291 5389 -11235
rect 5455 -11291 5691 -11235
rect -4159 -11399 5691 -11291
rect -4365 -11409 -4159 -11399
rect 5691 -11409 5897 -11399
<< via2 >>
rect 2408 1425 4098 1715
rect -2566 725 -876 1005
rect -2566 -589 -2222 -309
rect -2222 -589 -2164 -309
rect -2164 -589 -1750 -309
rect -1750 -589 -1692 -309
rect -1692 -589 -1278 -309
rect -1278 -589 -1220 -309
rect -1220 -589 -876 -309
rect -2668 -1289 -2576 -1009
rect -2576 -1289 -2518 -1009
rect -2518 -1289 -2340 -1009
rect -2340 -1289 -2282 -1009
rect -2282 -1289 -2104 -1009
rect -2104 -1289 -2046 -1009
rect -2046 -1289 -1868 -1009
rect -1868 -1289 -1810 -1009
rect -1810 -1289 -1632 -1009
rect -1632 -1289 -1574 -1009
rect -1574 -1289 -1396 -1009
rect -1396 -1289 -1338 -1009
rect -1338 -1289 -1160 -1009
rect -1160 -1289 -1102 -1009
rect -1102 -1289 -924 -1009
rect -924 -1289 -876 -1009
rect -50 -1080 5 -537
rect 5 -1080 263 -537
rect 263 -1080 321 -537
rect 321 -1080 394 -537
rect 1138 -1080 1211 -537
rect 1211 -1080 1269 -537
rect 1269 -1080 1527 -537
rect 1527 -1080 1582 -537
rect 2408 -589 2752 -309
rect 2752 -589 2810 -309
rect 2810 -589 3224 -309
rect 3224 -589 3282 -309
rect 3282 -589 3696 -309
rect 3696 -589 3754 -309
rect 3754 -589 4098 -309
rect 2409 -1289 2456 -1009
rect 2456 -1289 2634 -1009
rect 2634 -1289 2692 -1009
rect 2692 -1289 2870 -1009
rect 2870 -1289 2928 -1009
rect 2928 -1289 3106 -1009
rect 3106 -1289 3164 -1009
rect 3164 -1289 3342 -1009
rect 3342 -1289 3400 -1009
rect 3400 -1289 3578 -1009
rect 3578 -1289 3636 -1009
rect 3636 -1289 3814 -1009
rect 3814 -1289 3872 -1009
rect 3872 -1289 4050 -1009
rect 4050 -1289 4108 -1009
rect 4108 -1289 4201 -1009
rect -1132 -2948 -688 -2655
rect -50 -2948 394 -2655
rect 1138 -2948 1582 -2655
rect 2220 -2948 2664 -2655
rect -593 -3635 -553 -3342
rect -553 -3635 -495 -3342
rect -495 -3635 -149 -3342
rect 1677 -3635 2027 -3342
rect 2027 -3635 2085 -3342
rect 2085 -3635 2121 -3342
rect -1132 -4425 -688 -4272
rect -50 -4425 394 -4272
rect 1138 -4425 1582 -4272
rect 2220 -4425 2664 -4272
rect -593 -4679 -149 -4581
rect 1677 -4679 2121 -4581
rect -593 -4735 -467 -4679
rect -467 -4735 -401 -4679
rect -401 -4735 -275 -4679
rect -275 -4735 -209 -4679
rect -209 -4735 -149 -4679
rect 1677 -4735 1711 -4679
rect 1711 -4735 1837 -4679
rect 1837 -4735 1903 -4679
rect 1903 -4735 2029 -4679
rect 2029 -4735 2095 -4679
rect 2095 -4735 2121 -4679
<< metal3 >>
rect 2398 1715 4108 1725
rect -2576 1005 -866 1715
rect -2576 725 -2566 1005
rect -876 725 -866 1005
rect -2576 -309 -866 725
rect -2576 -589 -2566 -309
rect -876 -589 -866 -309
rect 2398 1425 2408 1715
rect 4098 1425 4108 1715
rect 2398 -309 4108 1425
rect -2576 -599 -866 -589
rect -60 -537 404 -527
rect -2678 -1009 -866 -1004
rect -2678 -1289 -2668 -1009
rect -876 -1289 -866 -1009
rect -2678 -1294 -866 -1289
rect -60 -1080 -50 -537
rect 394 -1080 404 -537
rect -1142 -2655 -678 -2645
rect -1142 -2948 -1132 -2655
rect -688 -2948 -678 -2655
rect -1142 -4272 -678 -2948
rect -60 -2655 404 -1080
rect -60 -2948 -50 -2655
rect 394 -2948 404 -2655
rect -1142 -4425 -1132 -4272
rect -688 -4425 -678 -4272
rect -1142 -4435 -678 -4425
rect -603 -3342 -139 -3332
rect -603 -3635 -593 -3342
rect -149 -3635 -139 -3342
rect -603 -4581 -139 -3635
rect -60 -4272 404 -2948
rect -60 -4425 -50 -4272
rect 394 -4425 404 -4272
rect -60 -4435 404 -4425
rect 1128 -537 1592 -527
rect 1128 -1080 1138 -537
rect 1582 -1080 1592 -537
rect 2398 -589 2408 -309
rect 4098 -589 4108 -309
rect 2398 -599 4108 -589
rect 1128 -2655 1592 -1080
rect 2399 -1009 4211 -1004
rect 2399 -1289 2409 -1009
rect 4201 -1289 4211 -1009
rect 2399 -1294 4211 -1289
rect 1128 -2948 1138 -2655
rect 1582 -2948 1592 -2655
rect 1128 -4272 1592 -2948
rect 2210 -2655 2674 -2645
rect 2210 -2948 2220 -2655
rect 2664 -2948 2674 -2655
rect 1128 -4425 1138 -4272
rect 1582 -4425 1592 -4272
rect 1128 -4435 1592 -4425
rect 1667 -3342 2131 -3332
rect 1667 -3635 1677 -3342
rect 2121 -3635 2131 -3342
rect -603 -4735 -593 -4581
rect -149 -4735 -139 -4581
rect -603 -4745 -139 -4735
rect 1667 -4581 2131 -3635
rect 2210 -4272 2674 -2948
rect 2210 -4425 2220 -4272
rect 2664 -4425 2674 -4272
rect 2210 -4435 2674 -4425
rect 1667 -4735 1677 -4581
rect 2121 -4735 2131 -4581
rect 1667 -4745 2131 -4735
<< via3 >>
rect -2668 -1289 -876 -1009
rect 2409 -1289 4201 -1009
<< metal4 >>
rect -4849 -1009 6381 -999
rect -4849 -1289 -2668 -1009
rect -876 -1289 2409 -1009
rect 4201 -1289 6381 -1009
rect -4849 -1299 6381 -1289
use sky130_fd_pr__nfet_01v8_2J7QF2  sky130_fd_pr__nfet_01v8_2J7QF2_0
timestamp 1697794388
transform 1 0 766 0 1 1215
box -737 -526 737 526
use sky130_fd_pr__nfet_01v8_U3DWQW  sky130_fd_pr__nfet_01v8_U3DWQW_0
timestamp 1697894789
transform 1 0 766 0 1 -799
box -819 -826 819 826
use sky130_fd_pr__nfet_01v8_Z85A38  sky130_fd_pr__nfet_01v8_Z85A38_0
timestamp 1697971722
transform 1 0 766 0 1 -3145
box -2351 -526 2351 526
use sky130_fd_pr__nfet_01v8_lvt_A3UXRA  sky130_fd_pr__nfet_01v8_lvt_A3UXRA_0
timestamp 1697808759
transform 1 0 766 0 1 -7985
box -4829 -3306 4829 3306
use sky130_fd_pr__pfet_01v8_477Z4B  sky130_fd_pr__pfet_01v8_477Z4B_0
timestamp 1698059623
transform 1 0 -1721 0 1 -799
box -993 -719 993 719
use sky130_fd_pr__pfet_01v8_477Z4B  sky130_fd_pr__pfet_01v8_477Z4B_1
timestamp 1698059623
transform 1 0 3253 0 1 -799
box -993 -719 993 719
<< labels >>
flabel metal2 6167 -3304 6472 -2986 0 FreeSans 1600 0 0 0 BIAS_CUR
port 6 nsew
flabel metal2 537 -3645 995 -3332 0 FreeSans 1600 0 0 0 VSS
flabel metal2 751 -4745 877 -4571 0 FreeSans 1600 0 0 0 VSS
flabel metal2 -4584 -4435 6208 -4262 0 FreeSans 1600 0 0 0 P1
flabel metal2 -237 -2958 737 -2645 0 FreeSans 1600 0 0 0 P1
flabel metal2 637 -1090 895 -527 0 FreeSans 1600 0 0 0 P1
flabel metal2 677 715 855 1015 0 FreeSans 1600 0 0 0 NEG2
flabel via1 737 1066 795 1366 0 FreeSans 1600 0 0 0 VSS
flabel metal2 -4849 -1985 -4544 -1667 0 FreeSans 1600 0 0 0 NEG
port 2 nsew
flabel metal2 479 -472 1053 8 0 FreeSans 1600 0 0 0 POS_D
flabel metal2 163 -1625 1369 -1145 0 FreeSans 1600 0 0 0 NEG_D
flabel metal2 -1928 -949 -1514 -649 0 FreeSans 1600 0 0 0 NEG_D
flabel via1 -1750 -599 -1692 -299 0 FreeSans 1600 0 0 0 NEG_2
flabel metal2 3046 -949 3460 -649 0 FreeSans 1600 0 0 0 POS_D
flabel metal2 3164 -1299 3342 -999 0 FreeSans 1600 0 0 0 VDD
flabel metal2 -1810 -1299 -1632 -999 0 FreeSans 1600 0 0 0 VDD
flabel metal2 -4849 1066 -4544 1379 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel via1 3224 -599 3282 -299 0 FreeSans 1600 0 0 0 EA_OUT
flabel metal2 29 1715 1503 2262 0 FreeSans 1600 0 0 0 EA_OUT
port 5 nsew
flabel metal4 -4849 -1299 -4544 -999 0 FreeSans 1600 0 0 0 VDD
port 4 nsew
flabel metal2 -4849 69 -4508 387 0 FreeSans 1600 0 0 0 POS
port 1 nsew
<< end >>
