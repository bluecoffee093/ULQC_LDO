magic
tech sky130A
magscale 1 2
timestamp 1697926267
<< nwell >>
rect -5457 -3219 5457 3219
<< pmoslvt >>
rect -5261 -3000 -4261 3000
rect -4203 -3000 -3203 3000
rect -3145 -3000 -2145 3000
rect -2087 -3000 -1087 3000
rect -1029 -3000 -29 3000
rect 29 -3000 1029 3000
rect 1087 -3000 2087 3000
rect 2145 -3000 3145 3000
rect 3203 -3000 4203 3000
rect 4261 -3000 5261 3000
<< pdiff >>
rect -5319 2988 -5261 3000
rect -5319 -2988 -5307 2988
rect -5273 -2988 -5261 2988
rect -5319 -3000 -5261 -2988
rect -4261 2988 -4203 3000
rect -4261 -2988 -4249 2988
rect -4215 -2988 -4203 2988
rect -4261 -3000 -4203 -2988
rect -3203 2988 -3145 3000
rect -3203 -2988 -3191 2988
rect -3157 -2988 -3145 2988
rect -3203 -3000 -3145 -2988
rect -2145 2988 -2087 3000
rect -2145 -2988 -2133 2988
rect -2099 -2988 -2087 2988
rect -2145 -3000 -2087 -2988
rect -1087 2988 -1029 3000
rect -1087 -2988 -1075 2988
rect -1041 -2988 -1029 2988
rect -1087 -3000 -1029 -2988
rect -29 2988 29 3000
rect -29 -2988 -17 2988
rect 17 -2988 29 2988
rect -29 -3000 29 -2988
rect 1029 2988 1087 3000
rect 1029 -2988 1041 2988
rect 1075 -2988 1087 2988
rect 1029 -3000 1087 -2988
rect 2087 2988 2145 3000
rect 2087 -2988 2099 2988
rect 2133 -2988 2145 2988
rect 2087 -3000 2145 -2988
rect 3145 2988 3203 3000
rect 3145 -2988 3157 2988
rect 3191 -2988 3203 2988
rect 3145 -3000 3203 -2988
rect 4203 2988 4261 3000
rect 4203 -2988 4215 2988
rect 4249 -2988 4261 2988
rect 4203 -3000 4261 -2988
rect 5261 2988 5319 3000
rect 5261 -2988 5273 2988
rect 5307 -2988 5319 2988
rect 5261 -3000 5319 -2988
<< pdiffc >>
rect -5307 -2988 -5273 2988
rect -4249 -2988 -4215 2988
rect -3191 -2988 -3157 2988
rect -2133 -2988 -2099 2988
rect -1075 -2988 -1041 2988
rect -17 -2988 17 2988
rect 1041 -2988 1075 2988
rect 2099 -2988 2133 2988
rect 3157 -2988 3191 2988
rect 4215 -2988 4249 2988
rect 5273 -2988 5307 2988
<< nsubdiff >>
rect -5421 3149 -5325 3183
rect 5325 3149 5421 3183
rect -5421 3087 -5387 3149
rect 5387 3087 5421 3149
rect -5421 -3149 -5387 -3087
rect 5387 -3149 5421 -3087
rect -5421 -3183 -5325 -3149
rect 5325 -3183 5421 -3149
<< nsubdiffcont >>
rect -5325 3149 5325 3183
rect -5421 -3087 -5387 3087
rect 5387 -3087 5421 3087
rect -5325 -3183 5325 -3149
<< poly >>
rect -5261 3081 -4261 3097
rect -5261 3047 -5245 3081
rect -4277 3047 -4261 3081
rect -5261 3000 -4261 3047
rect -4203 3081 -3203 3097
rect -4203 3047 -4187 3081
rect -3219 3047 -3203 3081
rect -4203 3000 -3203 3047
rect -3145 3081 -2145 3097
rect -3145 3047 -3129 3081
rect -2161 3047 -2145 3081
rect -3145 3000 -2145 3047
rect -2087 3081 -1087 3097
rect -2087 3047 -2071 3081
rect -1103 3047 -1087 3081
rect -2087 3000 -1087 3047
rect -1029 3081 -29 3097
rect -1029 3047 -1013 3081
rect -45 3047 -29 3081
rect -1029 3000 -29 3047
rect 29 3081 1029 3097
rect 29 3047 45 3081
rect 1013 3047 1029 3081
rect 29 3000 1029 3047
rect 1087 3081 2087 3097
rect 1087 3047 1103 3081
rect 2071 3047 2087 3081
rect 1087 3000 2087 3047
rect 2145 3081 3145 3097
rect 2145 3047 2161 3081
rect 3129 3047 3145 3081
rect 2145 3000 3145 3047
rect 3203 3081 4203 3097
rect 3203 3047 3219 3081
rect 4187 3047 4203 3081
rect 3203 3000 4203 3047
rect 4261 3081 5261 3097
rect 4261 3047 4277 3081
rect 5245 3047 5261 3081
rect 4261 3000 5261 3047
rect -5261 -3047 -4261 -3000
rect -5261 -3081 -5245 -3047
rect -4277 -3081 -4261 -3047
rect -5261 -3097 -4261 -3081
rect -4203 -3047 -3203 -3000
rect -4203 -3081 -4187 -3047
rect -3219 -3081 -3203 -3047
rect -4203 -3097 -3203 -3081
rect -3145 -3047 -2145 -3000
rect -3145 -3081 -3129 -3047
rect -2161 -3081 -2145 -3047
rect -3145 -3097 -2145 -3081
rect -2087 -3047 -1087 -3000
rect -2087 -3081 -2071 -3047
rect -1103 -3081 -1087 -3047
rect -2087 -3097 -1087 -3081
rect -1029 -3047 -29 -3000
rect -1029 -3081 -1013 -3047
rect -45 -3081 -29 -3047
rect -1029 -3097 -29 -3081
rect 29 -3047 1029 -3000
rect 29 -3081 45 -3047
rect 1013 -3081 1029 -3047
rect 29 -3097 1029 -3081
rect 1087 -3047 2087 -3000
rect 1087 -3081 1103 -3047
rect 2071 -3081 2087 -3047
rect 1087 -3097 2087 -3081
rect 2145 -3047 3145 -3000
rect 2145 -3081 2161 -3047
rect 3129 -3081 3145 -3047
rect 2145 -3097 3145 -3081
rect 3203 -3047 4203 -3000
rect 3203 -3081 3219 -3047
rect 4187 -3081 4203 -3047
rect 3203 -3097 4203 -3081
rect 4261 -3047 5261 -3000
rect 4261 -3081 4277 -3047
rect 5245 -3081 5261 -3047
rect 4261 -3097 5261 -3081
<< polycont >>
rect -5245 3047 -4277 3081
rect -4187 3047 -3219 3081
rect -3129 3047 -2161 3081
rect -2071 3047 -1103 3081
rect -1013 3047 -45 3081
rect 45 3047 1013 3081
rect 1103 3047 2071 3081
rect 2161 3047 3129 3081
rect 3219 3047 4187 3081
rect 4277 3047 5245 3081
rect -5245 -3081 -4277 -3047
rect -4187 -3081 -3219 -3047
rect -3129 -3081 -2161 -3047
rect -2071 -3081 -1103 -3047
rect -1013 -3081 -45 -3047
rect 45 -3081 1013 -3047
rect 1103 -3081 2071 -3047
rect 2161 -3081 3129 -3047
rect 3219 -3081 4187 -3047
rect 4277 -3081 5245 -3047
<< locali >>
rect -5421 3149 -5325 3183
rect 5325 3149 5421 3183
rect -5421 3087 -5387 3149
rect 5387 3087 5421 3149
rect -5261 3047 -5245 3081
rect -4277 3047 -4261 3081
rect -4203 3047 -4187 3081
rect -3219 3047 -3203 3081
rect -3145 3047 -3129 3081
rect -2161 3047 -2145 3081
rect -2087 3047 -2071 3081
rect -1103 3047 -1087 3081
rect -1029 3047 -1013 3081
rect -45 3047 -29 3081
rect 29 3047 45 3081
rect 1013 3047 1029 3081
rect 1087 3047 1103 3081
rect 2071 3047 2087 3081
rect 2145 3047 2161 3081
rect 3129 3047 3145 3081
rect 3203 3047 3219 3081
rect 4187 3047 4203 3081
rect 4261 3047 4277 3081
rect 5245 3047 5261 3081
rect -5307 2988 -5273 3004
rect -5307 -3004 -5273 -2988
rect -4249 2988 -4215 3004
rect -4249 -3004 -4215 -2988
rect -3191 2988 -3157 3004
rect -3191 -3004 -3157 -2988
rect -2133 2988 -2099 3004
rect -2133 -3004 -2099 -2988
rect -1075 2988 -1041 3004
rect -1075 -3004 -1041 -2988
rect -17 2988 17 3004
rect -17 -3004 17 -2988
rect 1041 2988 1075 3004
rect 1041 -3004 1075 -2988
rect 2099 2988 2133 3004
rect 2099 -3004 2133 -2988
rect 3157 2988 3191 3004
rect 3157 -3004 3191 -2988
rect 4215 2988 4249 3004
rect 4215 -3004 4249 -2988
rect 5273 2988 5307 3004
rect 5273 -3004 5307 -2988
rect -5261 -3081 -5245 -3047
rect -4277 -3081 -4261 -3047
rect -4203 -3081 -4187 -3047
rect -3219 -3081 -3203 -3047
rect -3145 -3081 -3129 -3047
rect -2161 -3081 -2145 -3047
rect -2087 -3081 -2071 -3047
rect -1103 -3081 -1087 -3047
rect -1029 -3081 -1013 -3047
rect -45 -3081 -29 -3047
rect 29 -3081 45 -3047
rect 1013 -3081 1029 -3047
rect 1087 -3081 1103 -3047
rect 2071 -3081 2087 -3047
rect 2145 -3081 2161 -3047
rect 3129 -3081 3145 -3047
rect 3203 -3081 3219 -3047
rect 4187 -3081 4203 -3047
rect 4261 -3081 4277 -3047
rect 5245 -3081 5261 -3047
rect -5421 -3149 -5387 -3087
rect 5387 -3149 5421 -3087
rect -5421 -3183 -5325 -3149
rect 5325 -3183 5421 -3149
<< viali >>
rect -5245 3047 -4277 3081
rect -4187 3047 -3219 3081
rect -3129 3047 -2161 3081
rect -2071 3047 -1103 3081
rect -1013 3047 -45 3081
rect 45 3047 1013 3081
rect 1103 3047 2071 3081
rect 2161 3047 3129 3081
rect 3219 3047 4187 3081
rect 4277 3047 5245 3081
rect -5307 -2988 -5273 2988
rect -4249 -2988 -4215 2988
rect -3191 -2988 -3157 2988
rect -2133 -2988 -2099 2988
rect -1075 -2988 -1041 2988
rect -17 -2988 17 2988
rect 1041 -2988 1075 2988
rect 2099 -2988 2133 2988
rect 3157 -2988 3191 2988
rect 4215 -2988 4249 2988
rect 5273 -2988 5307 2988
rect -5245 -3081 -4277 -3047
rect -4187 -3081 -3219 -3047
rect -3129 -3081 -2161 -3047
rect -2071 -3081 -1103 -3047
rect -1013 -3081 -45 -3047
rect 45 -3081 1013 -3047
rect 1103 -3081 2071 -3047
rect 2161 -3081 3129 -3047
rect 3219 -3081 4187 -3047
rect 4277 -3081 5245 -3047
<< metal1 >>
rect -5257 3081 -4265 3087
rect -5257 3047 -5245 3081
rect -4277 3047 -4265 3081
rect -5257 3041 -4265 3047
rect -4199 3081 -3207 3087
rect -4199 3047 -4187 3081
rect -3219 3047 -3207 3081
rect -4199 3041 -3207 3047
rect -3141 3081 -2149 3087
rect -3141 3047 -3129 3081
rect -2161 3047 -2149 3081
rect -3141 3041 -2149 3047
rect -2083 3081 -1091 3087
rect -2083 3047 -2071 3081
rect -1103 3047 -1091 3081
rect -2083 3041 -1091 3047
rect -1025 3081 -33 3087
rect -1025 3047 -1013 3081
rect -45 3047 -33 3081
rect -1025 3041 -33 3047
rect 33 3081 1025 3087
rect 33 3047 45 3081
rect 1013 3047 1025 3081
rect 33 3041 1025 3047
rect 1091 3081 2083 3087
rect 1091 3047 1103 3081
rect 2071 3047 2083 3081
rect 1091 3041 2083 3047
rect 2149 3081 3141 3087
rect 2149 3047 2161 3081
rect 3129 3047 3141 3081
rect 2149 3041 3141 3047
rect 3207 3081 4199 3087
rect 3207 3047 3219 3081
rect 4187 3047 4199 3081
rect 3207 3041 4199 3047
rect 4265 3081 5257 3087
rect 4265 3047 4277 3081
rect 5245 3047 5257 3081
rect 4265 3041 5257 3047
rect -5313 2988 -5267 3000
rect -5313 -2988 -5307 2988
rect -5273 -2988 -5267 2988
rect -5313 -3000 -5267 -2988
rect -4255 2988 -4209 3000
rect -4255 -2988 -4249 2988
rect -4215 -2988 -4209 2988
rect -4255 -3000 -4209 -2988
rect -3197 2988 -3151 3000
rect -3197 -2988 -3191 2988
rect -3157 -2988 -3151 2988
rect -3197 -3000 -3151 -2988
rect -2139 2988 -2093 3000
rect -2139 -2988 -2133 2988
rect -2099 -2988 -2093 2988
rect -2139 -3000 -2093 -2988
rect -1081 2988 -1035 3000
rect -1081 -2988 -1075 2988
rect -1041 -2988 -1035 2988
rect -1081 -3000 -1035 -2988
rect -23 2988 23 3000
rect -23 -2988 -17 2988
rect 17 -2988 23 2988
rect -23 -3000 23 -2988
rect 1035 2988 1081 3000
rect 1035 -2988 1041 2988
rect 1075 -2988 1081 2988
rect 1035 -3000 1081 -2988
rect 2093 2988 2139 3000
rect 2093 -2988 2099 2988
rect 2133 -2988 2139 2988
rect 2093 -3000 2139 -2988
rect 3151 2988 3197 3000
rect 3151 -2988 3157 2988
rect 3191 -2988 3197 2988
rect 3151 -3000 3197 -2988
rect 4209 2988 4255 3000
rect 4209 -2988 4215 2988
rect 4249 -2988 4255 2988
rect 4209 -3000 4255 -2988
rect 5267 2988 5313 3000
rect 5267 -2988 5273 2988
rect 5307 -2988 5313 2988
rect 5267 -3000 5313 -2988
rect -5257 -3047 -4265 -3041
rect -5257 -3081 -5245 -3047
rect -4277 -3081 -4265 -3047
rect -5257 -3087 -4265 -3081
rect -4199 -3047 -3207 -3041
rect -4199 -3081 -4187 -3047
rect -3219 -3081 -3207 -3047
rect -4199 -3087 -3207 -3081
rect -3141 -3047 -2149 -3041
rect -3141 -3081 -3129 -3047
rect -2161 -3081 -2149 -3047
rect -3141 -3087 -2149 -3081
rect -2083 -3047 -1091 -3041
rect -2083 -3081 -2071 -3047
rect -1103 -3081 -1091 -3047
rect -2083 -3087 -1091 -3081
rect -1025 -3047 -33 -3041
rect -1025 -3081 -1013 -3047
rect -45 -3081 -33 -3047
rect -1025 -3087 -33 -3081
rect 33 -3047 1025 -3041
rect 33 -3081 45 -3047
rect 1013 -3081 1025 -3047
rect 33 -3087 1025 -3081
rect 1091 -3047 2083 -3041
rect 1091 -3081 1103 -3047
rect 2071 -3081 2083 -3047
rect 1091 -3087 2083 -3081
rect 2149 -3047 3141 -3041
rect 2149 -3081 2161 -3047
rect 3129 -3081 3141 -3047
rect 2149 -3087 3141 -3081
rect 3207 -3047 4199 -3041
rect 3207 -3081 3219 -3047
rect 4187 -3081 4199 -3047
rect 3207 -3087 4199 -3081
rect 4265 -3047 5257 -3041
rect 4265 -3081 4277 -3047
rect 5245 -3081 5257 -3047
rect 4265 -3087 5257 -3081
<< properties >>
string FIXED_BBOX -5404 -3166 5404 3166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 30.0 l 5.0 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
