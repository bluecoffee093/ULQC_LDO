magic
tech sky130A
magscale 1 2
timestamp 1695858594
<< locali >>
rect 4277 -1001 4344 -931
rect 4701 -1000 4768 -929
rect 5123 -999 5190 -929
rect 2538 -1156 2770 -1154
rect 2672 -1346 2770 -1156
rect 3260 -1348 3262 -1152
rect 3350 -1348 3468 -1152
rect 2610 -1914 2772 -1912
rect 2700 -2110 2772 -1914
<< viali >>
rect 4276 -931 4345 -877
rect 4700 -929 4769 -875
rect 5122 -929 5191 -875
rect 2538 -1346 2672 -1156
rect 3262 -1348 3350 -1152
rect 2610 -2110 2700 -1914
<< metal1 >>
rect 2811 -845 3011 -645
rect 3514 -740 3714 -676
rect 4094 -717 5364 -700
rect 3514 -807 3950 -740
rect 2864 -964 2955 -845
rect 3514 -876 3714 -807
rect 2870 -1118 2950 -964
rect 3580 -1072 3644 -876
rect 2532 -1153 2678 -1144
rect 2532 -1154 2883 -1153
rect 2474 -1156 2883 -1154
rect 2474 -1346 2538 -1156
rect 2672 -1346 2883 -1156
rect 2474 -1350 2883 -1346
rect 2474 -1354 2678 -1350
rect 2532 -1358 2678 -1354
rect 2977 -1522 3006 -1150
rect 3256 -1152 3356 -1140
rect 3152 -1348 3262 -1152
rect 3350 -1153 3356 -1152
rect 3350 -1348 3585 -1153
rect 3152 -1350 3585 -1348
rect 3152 -1352 3356 -1350
rect 3256 -1360 3356 -1352
rect 3670 -1522 3699 -1148
rect 2808 -1722 3008 -1522
rect 3480 -1722 3699 -1522
rect 2604 -1906 2706 -1902
rect 2442 -1913 2706 -1906
rect 2442 -1914 2890 -1913
rect 2442 -2106 2610 -1914
rect 2604 -2110 2610 -2106
rect 2700 -2110 2890 -1914
rect 2604 -2122 2706 -2110
rect 2977 -2115 3006 -1722
rect 3326 -1914 3586 -1904
rect 3162 -2112 3586 -1914
rect 3162 -2114 3381 -2112
rect 3670 -2113 3699 -1722
rect 2866 -2342 2954 -2150
rect 3577 -2302 3644 -2148
rect 3854 -2302 3950 -807
rect 4092 -875 5364 -717
rect 4092 -877 4700 -875
rect 4092 -917 4276 -877
rect 4094 -927 4276 -917
rect 4264 -931 4276 -927
rect 4345 -927 4700 -877
rect 4345 -931 4357 -927
rect 4264 -937 4357 -931
rect 4688 -929 4700 -927
rect 4769 -927 5122 -875
rect 4769 -929 4781 -927
rect 4688 -935 4781 -929
rect 5110 -929 5122 -927
rect 5191 -927 5364 -875
rect 5191 -929 5203 -927
rect 5110 -935 5203 -929
rect 4278 -1046 4345 -937
rect 4701 -1045 4768 -935
rect 5123 -1043 5190 -935
rect 4278 -1070 4375 -1046
rect 4226 -1531 4255 -1147
rect 4340 -1354 4375 -1070
rect 4674 -1069 4768 -1045
rect 5097 -1068 5190 -1043
rect 4674 -1353 4709 -1069
rect 4060 -1731 4260 -1531
rect 4793 -1534 4822 -1146
rect 5097 -1351 5132 -1068
rect 5215 -1527 5244 -1146
rect 4226 -2112 4255 -1731
rect 4676 -1734 4876 -1534
rect 5113 -1727 5313 -1527
rect 4338 -2168 4373 -1904
rect 2810 -2542 3010 -2342
rect 3577 -2369 3950 -2302
rect 4284 -2324 4373 -2168
rect 4673 -2186 4708 -1903
rect 4793 -2111 4822 -1734
rect 5096 -2185 5131 -1903
rect 5215 -2111 5244 -1727
rect 4673 -2324 4769 -2186
rect 5096 -2324 5193 -2185
rect 3854 -2370 3950 -2369
rect 4104 -2542 5374 -2324
use sky130_fd_pr__nfet_01v8_64QSBY  XM1
timestamp 1695551012
transform 1 0 2912 0 1 -2042
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM2
timestamp 1695551012
transform 1 0 2911 0 1 -1216
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64QSBY  XM3
timestamp 1695551012
transform 1 0 3611 0 1 -2041
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM4
timestamp 1695551012
transform 1 0 3611 0 1 -1216
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64QSBY  XM5
timestamp 1695551012
transform 1 0 4312 0 1 -2039
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM6
timestamp 1695551012
transform 1 0 4313 0 1 -1216
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64QSBY  XM7
timestamp 1695551012
transform 1 0 4735 0 1 -2039
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM8
timestamp 1695551012
transform 1 0 4735 0 1 -1214
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64QSBY  sky130_fd_pr__nfet_01v8_64QSBY_0
timestamp 1695551012
transform 1 0 5158 0 1 -2038
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  sky130_fd_pr__pfet_01v8_MGS3BN_0
timestamp 1695551012
transform 1 0 5157 0 1 -1213
box -211 -284 211 284
<< labels >>
flabel metal1 4092 -917 4292 -717 0 FreeSans 256 0 0 0 VIN3
port 14 nsew
flabel metal1 3480 -1722 3680 -1522 0 FreeSans 256 0 0 0 VOUT2
port 11 nsew
flabel metal1 4060 -1731 4260 -1531 0 FreeSans 256 0 0 0 VOUT3
port 13 nsew
flabel metal1 5113 -1727 5313 -1527 0 FreeSans 256 0 0 0 BGR_OUT
port 4 nsew
flabel metal1 4676 -1734 4876 -1534 0 FreeSans 256 0 0 0 EA_OUT
port 6 nsew
flabel metal1 2474 -1354 2674 -1154 0 FreeSans 256 0 0 0 VIN1
port 10 nsew
flabel metal1 3152 -1352 3352 -1152 0 FreeSans 256 0 0 0 VIN2
port 12 nsew
flabel metal1 3514 -876 3714 -676 0 FreeSans 256 0 0 0 ADJ
port 1 nsew
flabel metal1 2811 -845 3011 -645 0 FreeSans 256 0 0 0 BGRT1
port 2 nsew
flabel metal1 2810 -2542 3010 -2342 0 FreeSans 256 0 0 0 BGRT2
port 3 nsew
flabel metal1 2808 -1722 3008 -1522 0 FreeSans 256 0 0 0 VOUT1
port 9 nsew
flabel metal1 2442 -2106 2642 -1906 0 FreeSans 240 0 0 0 VSS1
port 5 nsew
flabel metal1 3162 -2114 3381 -1914 0 FreeSans 240 0 0 0 VSS2
port 7 nsew
flabel metal1 4112 -2540 4331 -2340 0 FreeSans 240 0 0 0 VSS3
port 8 nsew
<< end >>
