magic
tech sky130A
magscale 1 2
timestamp 1697921066
<< error_p >>
rect -605 281 -547 287
rect -413 281 -355 287
rect -221 281 -163 287
rect -29 281 29 287
rect 163 281 221 287
rect 355 281 413 287
rect 547 281 605 287
rect -605 247 -593 281
rect -413 247 -401 281
rect -221 247 -209 281
rect -29 247 -17 281
rect 163 247 175 281
rect 355 247 367 281
rect 547 247 559 281
rect -605 241 -547 247
rect -413 241 -355 247
rect -221 241 -163 247
rect -29 241 29 247
rect 163 241 221 247
rect 355 241 413 247
rect 547 241 605 247
rect -701 -247 -643 -241
rect -509 -247 -451 -241
rect -317 -247 -259 -241
rect -125 -247 -67 -241
rect 67 -247 125 -241
rect 259 -247 317 -241
rect 451 -247 509 -241
rect 643 -247 701 -241
rect -701 -281 -689 -247
rect -509 -281 -497 -247
rect -317 -281 -305 -247
rect -125 -281 -113 -247
rect 67 -281 79 -247
rect 259 -281 271 -247
rect 451 -281 463 -247
rect 643 -281 655 -247
rect -701 -287 -643 -281
rect -509 -287 -451 -281
rect -317 -287 -259 -281
rect -125 -287 -67 -281
rect 67 -287 125 -281
rect 259 -287 317 -281
rect 451 -287 509 -281
rect 643 -287 701 -281
<< nwell >>
rect -689 262 689 300
rect -785 -300 785 262
<< pmos >>
rect -687 -200 -657 200
rect -591 -200 -561 200
rect -495 -200 -465 200
rect -399 -200 -369 200
rect -303 -200 -273 200
rect -207 -200 -177 200
rect -111 -200 -81 200
rect -15 -200 15 200
rect 81 -200 111 200
rect 177 -200 207 200
rect 273 -200 303 200
rect 369 -200 399 200
rect 465 -200 495 200
rect 561 -200 591 200
rect 657 -200 687 200
<< pdiff >>
rect -749 188 -687 200
rect -749 -188 -737 188
rect -703 -188 -687 188
rect -749 -200 -687 -188
rect -657 188 -591 200
rect -657 -188 -641 188
rect -607 -188 -591 188
rect -657 -200 -591 -188
rect -561 188 -495 200
rect -561 -188 -545 188
rect -511 -188 -495 188
rect -561 -200 -495 -188
rect -465 188 -399 200
rect -465 -188 -449 188
rect -415 -188 -399 188
rect -465 -200 -399 -188
rect -369 188 -303 200
rect -369 -188 -353 188
rect -319 -188 -303 188
rect -369 -200 -303 -188
rect -273 188 -207 200
rect -273 -188 -257 188
rect -223 -188 -207 188
rect -273 -200 -207 -188
rect -177 188 -111 200
rect -177 -188 -161 188
rect -127 -188 -111 188
rect -177 -200 -111 -188
rect -81 188 -15 200
rect -81 -188 -65 188
rect -31 -188 -15 188
rect -81 -200 -15 -188
rect 15 188 81 200
rect 15 -188 31 188
rect 65 -188 81 188
rect 15 -200 81 -188
rect 111 188 177 200
rect 111 -188 127 188
rect 161 -188 177 188
rect 111 -200 177 -188
rect 207 188 273 200
rect 207 -188 223 188
rect 257 -188 273 188
rect 207 -200 273 -188
rect 303 188 369 200
rect 303 -188 319 188
rect 353 -188 369 188
rect 303 -200 369 -188
rect 399 188 465 200
rect 399 -188 415 188
rect 449 -188 465 188
rect 399 -200 465 -188
rect 495 188 561 200
rect 495 -188 511 188
rect 545 -188 561 188
rect 495 -200 561 -188
rect 591 188 657 200
rect 591 -188 607 188
rect 641 -188 657 188
rect 591 -200 657 -188
rect 687 188 749 200
rect 687 -188 703 188
rect 737 -188 749 188
rect 687 -200 749 -188
<< pdiffc >>
rect -737 -188 -703 188
rect -641 -188 -607 188
rect -545 -188 -511 188
rect -449 -188 -415 188
rect -353 -188 -319 188
rect -257 -188 -223 188
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
rect 223 -188 257 188
rect 319 -188 353 188
rect 415 -188 449 188
rect 511 -188 545 188
rect 607 -188 641 188
rect 703 -188 737 188
<< poly >>
rect -609 281 -543 297
rect -609 247 -593 281
rect -559 247 -543 281
rect -609 231 -543 247
rect -417 281 -351 297
rect -417 247 -401 281
rect -367 247 -351 281
rect -417 231 -351 247
rect -225 281 -159 297
rect -225 247 -209 281
rect -175 247 -159 281
rect -225 231 -159 247
rect -33 281 33 297
rect -33 247 -17 281
rect 17 247 33 281
rect -33 231 33 247
rect 159 281 225 297
rect 159 247 175 281
rect 209 247 225 281
rect 159 231 225 247
rect 351 281 417 297
rect 351 247 367 281
rect 401 247 417 281
rect 351 231 417 247
rect 543 281 609 297
rect 543 247 559 281
rect 593 247 609 281
rect 543 231 609 247
rect -687 200 -657 226
rect -591 200 -561 231
rect -495 200 -465 226
rect -399 200 -369 231
rect -303 200 -273 226
rect -207 200 -177 231
rect -111 200 -81 226
rect -15 200 15 231
rect 81 200 111 226
rect 177 200 207 231
rect 273 200 303 226
rect 369 200 399 231
rect 465 200 495 226
rect 561 200 591 231
rect 657 200 687 226
rect -687 -231 -657 -200
rect -591 -226 -561 -200
rect -495 -231 -465 -200
rect -399 -226 -369 -200
rect -303 -231 -273 -200
rect -207 -226 -177 -200
rect -111 -231 -81 -200
rect -15 -226 15 -200
rect 81 -231 111 -200
rect 177 -226 207 -200
rect 273 -231 303 -200
rect 369 -226 399 -200
rect 465 -231 495 -200
rect 561 -226 591 -200
rect 657 -231 687 -200
rect -705 -247 -639 -231
rect -705 -281 -689 -247
rect -655 -281 -639 -247
rect -705 -297 -639 -281
rect -513 -247 -447 -231
rect -513 -281 -497 -247
rect -463 -281 -447 -247
rect -513 -297 -447 -281
rect -321 -247 -255 -231
rect -321 -281 -305 -247
rect -271 -281 -255 -247
rect -321 -297 -255 -281
rect -129 -247 -63 -231
rect -129 -281 -113 -247
rect -79 -281 -63 -247
rect -129 -297 -63 -281
rect 63 -247 129 -231
rect 63 -281 79 -247
rect 113 -281 129 -247
rect 63 -297 129 -281
rect 255 -247 321 -231
rect 255 -281 271 -247
rect 305 -281 321 -247
rect 255 -297 321 -281
rect 447 -247 513 -231
rect 447 -281 463 -247
rect 497 -281 513 -247
rect 447 -297 513 -281
rect 639 -247 705 -231
rect 639 -281 655 -247
rect 689 -281 705 -247
rect 639 -297 705 -281
<< polycont >>
rect -593 247 -559 281
rect -401 247 -367 281
rect -209 247 -175 281
rect -17 247 17 281
rect 175 247 209 281
rect 367 247 401 281
rect 559 247 593 281
rect -689 -281 -655 -247
rect -497 -281 -463 -247
rect -305 -281 -271 -247
rect -113 -281 -79 -247
rect 79 -281 113 -247
rect 271 -281 305 -247
rect 463 -281 497 -247
rect 655 -281 689 -247
<< locali >>
rect -609 247 -593 281
rect -559 247 -543 281
rect -417 247 -401 281
rect -367 247 -351 281
rect -225 247 -209 281
rect -175 247 -159 281
rect -33 247 -17 281
rect 17 247 33 281
rect 159 247 175 281
rect 209 247 225 281
rect 351 247 367 281
rect 401 247 417 281
rect 543 247 559 281
rect 593 247 609 281
rect -737 188 -703 204
rect -737 -204 -703 -188
rect -641 188 -607 204
rect -641 -204 -607 -188
rect -545 188 -511 204
rect -545 -204 -511 -188
rect -449 188 -415 204
rect -449 -204 -415 -188
rect -353 188 -319 204
rect -353 -204 -319 -188
rect -257 188 -223 204
rect -257 -204 -223 -188
rect -161 188 -127 204
rect -161 -204 -127 -188
rect -65 188 -31 204
rect -65 -204 -31 -188
rect 31 188 65 204
rect 31 -204 65 -188
rect 127 188 161 204
rect 127 -204 161 -188
rect 223 188 257 204
rect 223 -204 257 -188
rect 319 188 353 204
rect 319 -204 353 -188
rect 415 188 449 204
rect 415 -204 449 -188
rect 511 188 545 204
rect 511 -204 545 -188
rect 607 188 641 204
rect 607 -204 641 -188
rect 703 188 737 204
rect 703 -204 737 -188
rect -705 -281 -689 -247
rect -655 -281 -639 -247
rect -513 -281 -497 -247
rect -463 -281 -447 -247
rect -321 -281 -305 -247
rect -271 -281 -255 -247
rect -129 -281 -113 -247
rect -79 -281 -63 -247
rect 63 -281 79 -247
rect 113 -281 129 -247
rect 255 -281 271 -247
rect 305 -281 321 -247
rect 447 -281 463 -247
rect 497 -281 513 -247
rect 639 -281 655 -247
rect 689 -281 705 -247
<< viali >>
rect -593 247 -559 281
rect -401 247 -367 281
rect -209 247 -175 281
rect -17 247 17 281
rect 175 247 209 281
rect 367 247 401 281
rect 559 247 593 281
rect -737 -188 -703 188
rect -641 -188 -607 188
rect -545 -188 -511 188
rect -449 -188 -415 188
rect -353 -188 -319 188
rect -257 -188 -223 188
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
rect 223 -188 257 188
rect 319 -188 353 188
rect 415 -188 449 188
rect 511 -188 545 188
rect 607 -188 641 188
rect 703 -188 737 188
rect -689 -281 -655 -247
rect -497 -281 -463 -247
rect -305 -281 -271 -247
rect -113 -281 -79 -247
rect 79 -281 113 -247
rect 271 -281 305 -247
rect 463 -281 497 -247
rect 655 -281 689 -247
<< metal1 >>
rect -605 281 -547 287
rect -605 247 -593 281
rect -559 247 -547 281
rect -605 241 -547 247
rect -413 281 -355 287
rect -413 247 -401 281
rect -367 247 -355 281
rect -413 241 -355 247
rect -221 281 -163 287
rect -221 247 -209 281
rect -175 247 -163 281
rect -221 241 -163 247
rect -29 281 29 287
rect -29 247 -17 281
rect 17 247 29 281
rect -29 241 29 247
rect 163 281 221 287
rect 163 247 175 281
rect 209 247 221 281
rect 163 241 221 247
rect 355 281 413 287
rect 355 247 367 281
rect 401 247 413 281
rect 355 241 413 247
rect 547 281 605 287
rect 547 247 559 281
rect 593 247 605 281
rect 547 241 605 247
rect -743 188 -697 200
rect -743 -188 -737 188
rect -703 -188 -697 188
rect -743 -200 -697 -188
rect -647 188 -601 200
rect -647 -188 -641 188
rect -607 -188 -601 188
rect -647 -200 -601 -188
rect -551 188 -505 200
rect -551 -188 -545 188
rect -511 -188 -505 188
rect -551 -200 -505 -188
rect -455 188 -409 200
rect -455 -188 -449 188
rect -415 -188 -409 188
rect -455 -200 -409 -188
rect -359 188 -313 200
rect -359 -188 -353 188
rect -319 -188 -313 188
rect -359 -200 -313 -188
rect -263 188 -217 200
rect -263 -188 -257 188
rect -223 -188 -217 188
rect -263 -200 -217 -188
rect -167 188 -121 200
rect -167 -188 -161 188
rect -127 -188 -121 188
rect -167 -200 -121 -188
rect -71 188 -25 200
rect -71 -188 -65 188
rect -31 -188 -25 188
rect -71 -200 -25 -188
rect 25 188 71 200
rect 25 -188 31 188
rect 65 -188 71 188
rect 25 -200 71 -188
rect 121 188 167 200
rect 121 -188 127 188
rect 161 -188 167 188
rect 121 -200 167 -188
rect 217 188 263 200
rect 217 -188 223 188
rect 257 -188 263 188
rect 217 -200 263 -188
rect 313 188 359 200
rect 313 -188 319 188
rect 353 -188 359 188
rect 313 -200 359 -188
rect 409 188 455 200
rect 409 -188 415 188
rect 449 -188 455 188
rect 409 -200 455 -188
rect 505 188 551 200
rect 505 -188 511 188
rect 545 -188 551 188
rect 505 -200 551 -188
rect 601 188 647 200
rect 601 -188 607 188
rect 641 -188 647 188
rect 601 -200 647 -188
rect 697 188 743 200
rect 697 -188 703 188
rect 737 -188 743 188
rect 697 -200 743 -188
rect -701 -247 -643 -241
rect -701 -281 -689 -247
rect -655 -281 -643 -247
rect -701 -287 -643 -281
rect -509 -247 -451 -241
rect -509 -281 -497 -247
rect -463 -281 -451 -247
rect -509 -287 -451 -281
rect -317 -247 -259 -241
rect -317 -281 -305 -247
rect -271 -281 -259 -247
rect -317 -287 -259 -281
rect -125 -247 -67 -241
rect -125 -281 -113 -247
rect -79 -281 -67 -247
rect -125 -287 -67 -281
rect 67 -247 125 -241
rect 67 -281 79 -247
rect 113 -281 125 -247
rect 67 -287 125 -281
rect 259 -247 317 -241
rect 259 -281 271 -247
rect 305 -281 317 -247
rect 259 -287 317 -281
rect 451 -247 509 -241
rect 451 -281 463 -247
rect 497 -281 509 -247
rect 451 -287 509 -281
rect 643 -247 701 -241
rect 643 -281 655 -247
rect 689 -281 701 -247
rect 643 -287 701 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 1 nf 15 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
