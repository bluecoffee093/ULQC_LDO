magic
tech sky130A
timestamp 1697794388
<< error_p >>
rect -625 286 -596 289
rect -403 286 -374 289
rect -181 286 -152 289
rect 41 286 70 289
rect 263 286 292 289
rect 485 286 514 289
rect 707 286 736 289
rect -625 269 -619 286
rect -403 269 -397 286
rect -181 269 -175 286
rect 41 269 47 286
rect 263 269 269 286
rect 485 269 491 286
rect 707 269 713 286
rect -625 266 -596 269
rect -403 266 -374 269
rect -181 266 -152 269
rect 41 266 70 269
rect 263 266 292 269
rect 485 266 514 269
rect 707 266 736 269
rect -736 -269 -707 -266
rect -514 -269 -485 -266
rect -292 -269 -263 -266
rect -70 -269 -41 -266
rect 152 -269 181 -266
rect 374 -269 403 -266
rect 596 -269 625 -266
rect -736 -286 -730 -269
rect -514 -286 -508 -269
rect -292 -286 -286 -269
rect -70 -286 -64 -269
rect 152 -286 158 -269
rect 374 -286 380 -269
rect 596 -286 602 -269
rect -736 -289 -707 -286
rect -514 -289 -485 -286
rect -292 -289 -263 -286
rect -70 -289 -41 -286
rect 152 -289 181 -286
rect 374 -289 403 -286
rect 596 -289 625 -286
<< nmos >>
rect -734 -250 -709 250
rect -623 -250 -598 250
rect -512 -250 -487 250
rect -401 -250 -376 250
rect -290 -250 -265 250
rect -179 -250 -154 250
rect -68 -250 -43 250
rect 43 -250 68 250
rect 154 -250 179 250
rect 265 -250 290 250
rect 376 -250 401 250
rect 487 -250 512 250
rect 598 -250 623 250
rect 709 -250 734 250
<< ndiff >>
rect -763 244 -734 250
rect -763 -244 -757 244
rect -740 -244 -734 244
rect -763 -250 -734 -244
rect -709 244 -680 250
rect -709 -244 -703 244
rect -686 -244 -680 244
rect -709 -250 -680 -244
rect -652 244 -623 250
rect -652 -244 -646 244
rect -629 -244 -623 244
rect -652 -250 -623 -244
rect -598 244 -569 250
rect -598 -244 -592 244
rect -575 -244 -569 244
rect -598 -250 -569 -244
rect -541 244 -512 250
rect -541 -244 -535 244
rect -518 -244 -512 244
rect -541 -250 -512 -244
rect -487 244 -458 250
rect -487 -244 -481 244
rect -464 -244 -458 244
rect -487 -250 -458 -244
rect -430 244 -401 250
rect -430 -244 -424 244
rect -407 -244 -401 244
rect -430 -250 -401 -244
rect -376 244 -347 250
rect -376 -244 -370 244
rect -353 -244 -347 244
rect -376 -250 -347 -244
rect -319 244 -290 250
rect -319 -244 -313 244
rect -296 -244 -290 244
rect -319 -250 -290 -244
rect -265 244 -236 250
rect -265 -244 -259 244
rect -242 -244 -236 244
rect -265 -250 -236 -244
rect -208 244 -179 250
rect -208 -244 -202 244
rect -185 -244 -179 244
rect -208 -250 -179 -244
rect -154 244 -125 250
rect -154 -244 -148 244
rect -131 -244 -125 244
rect -154 -250 -125 -244
rect -97 244 -68 250
rect -97 -244 -91 244
rect -74 -244 -68 244
rect -97 -250 -68 -244
rect -43 244 -14 250
rect -43 -244 -37 244
rect -20 -244 -14 244
rect -43 -250 -14 -244
rect 14 244 43 250
rect 14 -244 20 244
rect 37 -244 43 244
rect 14 -250 43 -244
rect 68 244 97 250
rect 68 -244 74 244
rect 91 -244 97 244
rect 68 -250 97 -244
rect 125 244 154 250
rect 125 -244 131 244
rect 148 -244 154 244
rect 125 -250 154 -244
rect 179 244 208 250
rect 179 -244 185 244
rect 202 -244 208 244
rect 179 -250 208 -244
rect 236 244 265 250
rect 236 -244 242 244
rect 259 -244 265 244
rect 236 -250 265 -244
rect 290 244 319 250
rect 290 -244 296 244
rect 313 -244 319 244
rect 290 -250 319 -244
rect 347 244 376 250
rect 347 -244 353 244
rect 370 -244 376 244
rect 347 -250 376 -244
rect 401 244 430 250
rect 401 -244 407 244
rect 424 -244 430 244
rect 401 -250 430 -244
rect 458 244 487 250
rect 458 -244 464 244
rect 481 -244 487 244
rect 458 -250 487 -244
rect 512 244 541 250
rect 512 -244 518 244
rect 535 -244 541 244
rect 512 -250 541 -244
rect 569 244 598 250
rect 569 -244 575 244
rect 592 -244 598 244
rect 569 -250 598 -244
rect 623 244 652 250
rect 623 -244 629 244
rect 646 -244 652 244
rect 623 -250 652 -244
rect 680 244 709 250
rect 680 -244 686 244
rect 703 -244 709 244
rect 680 -250 709 -244
rect 734 244 763 250
rect 734 -244 740 244
rect 757 -244 763 244
rect 734 -250 763 -244
<< ndiffc >>
rect -757 -244 -740 244
rect -703 -244 -686 244
rect -646 -244 -629 244
rect -592 -244 -575 244
rect -535 -244 -518 244
rect -481 -244 -464 244
rect -424 -244 -407 244
rect -370 -244 -353 244
rect -313 -244 -296 244
rect -259 -244 -242 244
rect -202 -244 -185 244
rect -148 -244 -131 244
rect -91 -244 -74 244
rect -37 -244 -20 244
rect 20 -244 37 244
rect 74 -244 91 244
rect 131 -244 148 244
rect 185 -244 202 244
rect 242 -244 259 244
rect 296 -244 313 244
rect 353 -244 370 244
rect 407 -244 424 244
rect 464 -244 481 244
rect 518 -244 535 244
rect 575 -244 592 244
rect 629 -244 646 244
rect 686 -244 703 244
rect 740 -244 757 244
<< poly >>
rect -627 286 -594 294
rect -627 269 -619 286
rect -602 269 -594 286
rect -734 250 -709 263
rect -627 261 -594 269
rect -405 286 -372 294
rect -405 269 -397 286
rect -380 269 -372 286
rect -623 250 -598 261
rect -512 250 -487 263
rect -405 261 -372 269
rect -183 286 -150 294
rect -183 269 -175 286
rect -158 269 -150 286
rect -401 250 -376 261
rect -290 250 -265 263
rect -183 261 -150 269
rect 39 286 72 294
rect 39 269 47 286
rect 64 269 72 286
rect -179 250 -154 261
rect -68 250 -43 263
rect 39 261 72 269
rect 261 286 294 294
rect 261 269 269 286
rect 286 269 294 286
rect 43 250 68 261
rect 154 250 179 263
rect 261 261 294 269
rect 483 286 516 294
rect 483 269 491 286
rect 508 269 516 286
rect 265 250 290 261
rect 376 250 401 263
rect 483 261 516 269
rect 705 286 738 294
rect 705 269 713 286
rect 730 269 738 286
rect 487 250 512 261
rect 598 250 623 263
rect 705 261 738 269
rect 709 250 734 261
rect -734 -261 -709 -250
rect -738 -269 -705 -261
rect -623 -263 -598 -250
rect -512 -261 -487 -250
rect -738 -286 -730 -269
rect -713 -286 -705 -269
rect -738 -294 -705 -286
rect -516 -269 -483 -261
rect -401 -263 -376 -250
rect -290 -261 -265 -250
rect -516 -286 -508 -269
rect -491 -286 -483 -269
rect -516 -294 -483 -286
rect -294 -269 -261 -261
rect -179 -263 -154 -250
rect -68 -261 -43 -250
rect -294 -286 -286 -269
rect -269 -286 -261 -269
rect -294 -294 -261 -286
rect -72 -269 -39 -261
rect 43 -263 68 -250
rect 154 -261 179 -250
rect -72 -286 -64 -269
rect -47 -286 -39 -269
rect -72 -294 -39 -286
rect 150 -269 183 -261
rect 265 -263 290 -250
rect 376 -261 401 -250
rect 150 -286 158 -269
rect 175 -286 183 -269
rect 150 -294 183 -286
rect 372 -269 405 -261
rect 487 -263 512 -250
rect 598 -261 623 -250
rect 372 -286 380 -269
rect 397 -286 405 -269
rect 372 -294 405 -286
rect 594 -269 627 -261
rect 709 -263 734 -250
rect 594 -286 602 -269
rect 619 -286 627 -269
rect 594 -294 627 -286
<< polycont >>
rect -619 269 -602 286
rect -397 269 -380 286
rect -175 269 -158 286
rect 47 269 64 286
rect 269 269 286 286
rect 491 269 508 286
rect 713 269 730 286
rect -730 -286 -713 -269
rect -508 -286 -491 -269
rect -286 -286 -269 -269
rect -64 -286 -47 -269
rect 158 -286 175 -269
rect 380 -286 397 -269
rect 602 -286 619 -269
<< locali >>
rect -627 269 -619 286
rect -602 269 -594 286
rect -405 269 -397 286
rect -380 269 -372 286
rect -183 269 -175 286
rect -158 269 -150 286
rect 39 269 47 286
rect 64 269 72 286
rect 261 269 269 286
rect 286 269 294 286
rect 483 269 491 286
rect 508 269 516 286
rect 705 269 713 286
rect 730 269 738 286
rect -757 244 -740 252
rect -757 -252 -740 -244
rect -703 244 -686 252
rect -703 -252 -686 -244
rect -646 244 -629 252
rect -646 -252 -629 -244
rect -592 244 -575 252
rect -592 -252 -575 -244
rect -535 244 -518 252
rect -535 -252 -518 -244
rect -481 244 -464 252
rect -481 -252 -464 -244
rect -424 244 -407 252
rect -424 -252 -407 -244
rect -370 244 -353 252
rect -370 -252 -353 -244
rect -313 244 -296 252
rect -313 -252 -296 -244
rect -259 244 -242 252
rect -259 -252 -242 -244
rect -202 244 -185 252
rect -202 -252 -185 -244
rect -148 244 -131 252
rect -148 -252 -131 -244
rect -91 244 -74 252
rect -91 -252 -74 -244
rect -37 244 -20 252
rect -37 -252 -20 -244
rect 20 244 37 252
rect 20 -252 37 -244
rect 74 244 91 252
rect 74 -252 91 -244
rect 131 244 148 252
rect 131 -252 148 -244
rect 185 244 202 252
rect 185 -252 202 -244
rect 242 244 259 252
rect 242 -252 259 -244
rect 296 244 313 252
rect 296 -252 313 -244
rect 353 244 370 252
rect 353 -252 370 -244
rect 407 244 424 252
rect 407 -252 424 -244
rect 464 244 481 252
rect 464 -252 481 -244
rect 518 244 535 252
rect 518 -252 535 -244
rect 575 244 592 252
rect 575 -252 592 -244
rect 629 244 646 252
rect 629 -252 646 -244
rect 686 244 703 252
rect 686 -252 703 -244
rect 740 244 757 252
rect 740 -252 757 -244
rect -738 -286 -730 -269
rect -713 -286 -705 -269
rect -516 -286 -508 -269
rect -491 -286 -483 -269
rect -294 -286 -286 -269
rect -269 -286 -261 -269
rect -72 -286 -64 -269
rect -47 -286 -39 -269
rect 150 -286 158 -269
rect 175 -286 183 -269
rect 372 -286 380 -269
rect 397 -286 405 -269
rect 594 -286 602 -269
rect 619 -286 627 -269
<< viali >>
rect -619 269 -602 286
rect -397 269 -380 286
rect -175 269 -158 286
rect 47 269 64 286
rect 269 269 286 286
rect 491 269 508 286
rect 713 269 730 286
rect -757 -244 -740 244
rect -703 -244 -686 244
rect -646 -244 -629 244
rect -592 -244 -575 244
rect -535 -244 -518 244
rect -481 -244 -464 244
rect -424 -244 -407 244
rect -370 -244 -353 244
rect -313 -244 -296 244
rect -259 -244 -242 244
rect -202 -244 -185 244
rect -148 -244 -131 244
rect -91 -244 -74 244
rect -37 -244 -20 244
rect 20 -244 37 244
rect 74 -244 91 244
rect 131 -244 148 244
rect 185 -244 202 244
rect 242 -244 259 244
rect 296 -244 313 244
rect 353 -244 370 244
rect 407 -244 424 244
rect 464 -244 481 244
rect 518 -244 535 244
rect 575 -244 592 244
rect 629 -244 646 244
rect 686 -244 703 244
rect 740 -244 757 244
rect -730 -286 -713 -269
rect -508 -286 -491 -269
rect -286 -286 -269 -269
rect -64 -286 -47 -269
rect 158 -286 175 -269
rect 380 -286 397 -269
rect 602 -286 619 -269
<< metal1 >>
rect -625 286 -596 289
rect -625 269 -619 286
rect -602 269 -596 286
rect -625 266 -596 269
rect -403 286 -374 289
rect -403 269 -397 286
rect -380 269 -374 286
rect -403 266 -374 269
rect -181 286 -152 289
rect -181 269 -175 286
rect -158 269 -152 286
rect -181 266 -152 269
rect 41 286 70 289
rect 41 269 47 286
rect 64 269 70 286
rect 41 266 70 269
rect 263 286 292 289
rect 263 269 269 286
rect 286 269 292 286
rect 263 266 292 269
rect 485 286 514 289
rect 485 269 491 286
rect 508 269 514 286
rect 485 266 514 269
rect 707 286 736 289
rect 707 269 713 286
rect 730 269 736 286
rect 707 266 736 269
rect -760 244 -737 250
rect -760 -244 -757 244
rect -740 -244 -737 244
rect -760 -250 -737 -244
rect -706 244 -683 250
rect -706 -244 -703 244
rect -686 -244 -683 244
rect -706 -250 -683 -244
rect -649 244 -626 250
rect -649 -244 -646 244
rect -629 -244 -626 244
rect -649 -250 -626 -244
rect -595 244 -572 250
rect -595 -244 -592 244
rect -575 -244 -572 244
rect -595 -250 -572 -244
rect -538 244 -515 250
rect -538 -244 -535 244
rect -518 -244 -515 244
rect -538 -250 -515 -244
rect -484 244 -461 250
rect -484 -244 -481 244
rect -464 -244 -461 244
rect -484 -250 -461 -244
rect -427 244 -404 250
rect -427 -244 -424 244
rect -407 -244 -404 244
rect -427 -250 -404 -244
rect -373 244 -350 250
rect -373 -244 -370 244
rect -353 -244 -350 244
rect -373 -250 -350 -244
rect -316 244 -293 250
rect -316 -244 -313 244
rect -296 -244 -293 244
rect -316 -250 -293 -244
rect -262 244 -239 250
rect -262 -244 -259 244
rect -242 -244 -239 244
rect -262 -250 -239 -244
rect -205 244 -182 250
rect -205 -244 -202 244
rect -185 -244 -182 244
rect -205 -250 -182 -244
rect -151 244 -128 250
rect -151 -244 -148 244
rect -131 -244 -128 244
rect -151 -250 -128 -244
rect -94 244 -71 250
rect -94 -244 -91 244
rect -74 -244 -71 244
rect -94 -250 -71 -244
rect -40 244 -17 250
rect -40 -244 -37 244
rect -20 -244 -17 244
rect -40 -250 -17 -244
rect 17 244 40 250
rect 17 -244 20 244
rect 37 -244 40 244
rect 17 -250 40 -244
rect 71 244 94 250
rect 71 -244 74 244
rect 91 -244 94 244
rect 71 -250 94 -244
rect 128 244 151 250
rect 128 -244 131 244
rect 148 -244 151 244
rect 128 -250 151 -244
rect 182 244 205 250
rect 182 -244 185 244
rect 202 -244 205 244
rect 182 -250 205 -244
rect 239 244 262 250
rect 239 -244 242 244
rect 259 -244 262 244
rect 239 -250 262 -244
rect 293 244 316 250
rect 293 -244 296 244
rect 313 -244 316 244
rect 293 -250 316 -244
rect 350 244 373 250
rect 350 -244 353 244
rect 370 -244 373 244
rect 350 -250 373 -244
rect 404 244 427 250
rect 404 -244 407 244
rect 424 -244 427 244
rect 404 -250 427 -244
rect 461 244 484 250
rect 461 -244 464 244
rect 481 -244 484 244
rect 461 -250 484 -244
rect 515 244 538 250
rect 515 -244 518 244
rect 535 -244 538 244
rect 515 -250 538 -244
rect 572 244 595 250
rect 572 -244 575 244
rect 592 -244 595 244
rect 572 -250 595 -244
rect 626 244 649 250
rect 626 -244 629 244
rect 646 -244 649 244
rect 626 -250 649 -244
rect 683 244 706 250
rect 683 -244 686 244
rect 703 -244 706 244
rect 683 -250 706 -244
rect 737 244 760 250
rect 737 -244 740 244
rect 757 -244 760 244
rect 737 -250 760 -244
rect -736 -269 -707 -266
rect -736 -286 -730 -269
rect -713 -286 -707 -269
rect -736 -289 -707 -286
rect -514 -269 -485 -266
rect -514 -286 -508 -269
rect -491 -286 -485 -269
rect -514 -289 -485 -286
rect -292 -269 -263 -266
rect -292 -286 -286 -269
rect -269 -286 -263 -269
rect -292 -289 -263 -286
rect -70 -269 -41 -266
rect -70 -286 -64 -269
rect -47 -286 -41 -269
rect -70 -289 -41 -286
rect 152 -269 181 -266
rect 152 -286 158 -269
rect 175 -286 181 -269
rect 152 -289 181 -286
rect 374 -269 403 -266
rect 374 -286 380 -269
rect 397 -286 403 -269
rect 374 -289 403 -286
rect 596 -269 625 -266
rect 596 -286 602 -269
rect 619 -286 625 -269
rect 596 -289 625 -286
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.25 m 1 nf 14 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
