** sch_path: /foss/designs/ulqc_ldo/repo/ULQC_LDO/xschem/bandgap.sch
**.subckt bandgap
XM4 vg_n vg_n v1 VSS sky130_fd_pr__nfet_01v8 L=10 W=60 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
XQ1 VSS VSS net2 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
V1 VDD VSS 1.8
.save i(v1)
XQ3 VSS VSS net3 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
R1 Vout v_iptat 250k m=1
XQ2 VSS VSS v3 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=8
R2 net1 v3 28k m=1
V2 VSS GND 0
.save i(v2)
Vmeas1 v1 net2 0
.save i(vmeas1)
Vmeas2 v2 net1 0
.save i(vmeas2)
Vmeas3 v_iptat net3 0
.save i(vmeas3)
XM1 vg_n vg_p VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=60 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
XM2 vg_p vg_p VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=60 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
XM3 vg_p vg_n v2 VSS sky130_fd_pr__nfet_01v8 L=10 W=60 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
XM5 Vout vg_p VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=60 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
**** begin user architecture code


* ngspice commands
.control
save all
save @m.xm1.msky130_fd_pr__pfet_01v8_lvt[vth]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[vth]
*dc temp -40 125 0.1
dc V1 1.2 2.5 0.01
plot v(Vout)
*op
write bandgap.raw
.endc



**** end user architecture code
.end
