magic
tech sky130A
magscale 1 2
timestamp 1697815432
<< nmos >>
rect -2293 47 -2093 547
rect -2035 47 -1835 547
rect -1777 47 -1577 547
rect -1519 47 -1319 547
rect -1261 47 -1061 547
rect -1003 47 -803 547
rect -745 47 -545 547
rect -487 47 -287 547
rect -229 47 -29 547
rect 29 47 229 547
rect 287 47 487 547
rect 545 47 745 547
rect 803 47 1003 547
rect 1061 47 1261 547
rect 1319 47 1519 547
rect 1577 47 1777 547
rect 1835 47 2035 547
rect 2093 47 2293 547
rect -2293 -547 -2093 -47
rect -2035 -547 -1835 -47
rect -1777 -547 -1577 -47
rect -1519 -547 -1319 -47
rect -1261 -547 -1061 -47
rect -1003 -547 -803 -47
rect -745 -547 -545 -47
rect -487 -547 -287 -47
rect -229 -547 -29 -47
rect 29 -547 229 -47
rect 287 -547 487 -47
rect 545 -547 745 -47
rect 803 -547 1003 -47
rect 1061 -547 1261 -47
rect 1319 -547 1519 -47
rect 1577 -547 1777 -47
rect 1835 -547 2035 -47
rect 2093 -547 2293 -47
<< ndiff >>
rect -2351 535 -2293 547
rect -2351 59 -2339 535
rect -2305 59 -2293 535
rect -2351 47 -2293 59
rect -2093 535 -2035 547
rect -2093 59 -2081 535
rect -2047 59 -2035 535
rect -2093 47 -2035 59
rect -1835 535 -1777 547
rect -1835 59 -1823 535
rect -1789 59 -1777 535
rect -1835 47 -1777 59
rect -1577 535 -1519 547
rect -1577 59 -1565 535
rect -1531 59 -1519 535
rect -1577 47 -1519 59
rect -1319 535 -1261 547
rect -1319 59 -1307 535
rect -1273 59 -1261 535
rect -1319 47 -1261 59
rect -1061 535 -1003 547
rect -1061 59 -1049 535
rect -1015 59 -1003 535
rect -1061 47 -1003 59
rect -803 535 -745 547
rect -803 59 -791 535
rect -757 59 -745 535
rect -803 47 -745 59
rect -545 535 -487 547
rect -545 59 -533 535
rect -499 59 -487 535
rect -545 47 -487 59
rect -287 535 -229 547
rect -287 59 -275 535
rect -241 59 -229 535
rect -287 47 -229 59
rect -29 535 29 547
rect -29 59 -17 535
rect 17 59 29 535
rect -29 47 29 59
rect 229 535 287 547
rect 229 59 241 535
rect 275 59 287 535
rect 229 47 287 59
rect 487 535 545 547
rect 487 59 499 535
rect 533 59 545 535
rect 487 47 545 59
rect 745 535 803 547
rect 745 59 757 535
rect 791 59 803 535
rect 745 47 803 59
rect 1003 535 1061 547
rect 1003 59 1015 535
rect 1049 59 1061 535
rect 1003 47 1061 59
rect 1261 535 1319 547
rect 1261 59 1273 535
rect 1307 59 1319 535
rect 1261 47 1319 59
rect 1519 535 1577 547
rect 1519 59 1531 535
rect 1565 59 1577 535
rect 1519 47 1577 59
rect 1777 535 1835 547
rect 1777 59 1789 535
rect 1823 59 1835 535
rect 1777 47 1835 59
rect 2035 535 2093 547
rect 2035 59 2047 535
rect 2081 59 2093 535
rect 2035 47 2093 59
rect 2293 535 2351 547
rect 2293 59 2305 535
rect 2339 59 2351 535
rect 2293 47 2351 59
rect -2351 -59 -2293 -47
rect -2351 -535 -2339 -59
rect -2305 -535 -2293 -59
rect -2351 -547 -2293 -535
rect -2093 -59 -2035 -47
rect -2093 -535 -2081 -59
rect -2047 -535 -2035 -59
rect -2093 -547 -2035 -535
rect -1835 -59 -1777 -47
rect -1835 -535 -1823 -59
rect -1789 -535 -1777 -59
rect -1835 -547 -1777 -535
rect -1577 -59 -1519 -47
rect -1577 -535 -1565 -59
rect -1531 -535 -1519 -59
rect -1577 -547 -1519 -535
rect -1319 -59 -1261 -47
rect -1319 -535 -1307 -59
rect -1273 -535 -1261 -59
rect -1319 -547 -1261 -535
rect -1061 -59 -1003 -47
rect -1061 -535 -1049 -59
rect -1015 -535 -1003 -59
rect -1061 -547 -1003 -535
rect -803 -59 -745 -47
rect -803 -535 -791 -59
rect -757 -535 -745 -59
rect -803 -547 -745 -535
rect -545 -59 -487 -47
rect -545 -535 -533 -59
rect -499 -535 -487 -59
rect -545 -547 -487 -535
rect -287 -59 -229 -47
rect -287 -535 -275 -59
rect -241 -535 -229 -59
rect -287 -547 -229 -535
rect -29 -59 29 -47
rect -29 -535 -17 -59
rect 17 -535 29 -59
rect -29 -547 29 -535
rect 229 -59 287 -47
rect 229 -535 241 -59
rect 275 -535 287 -59
rect 229 -547 287 -535
rect 487 -59 545 -47
rect 487 -535 499 -59
rect 533 -535 545 -59
rect 487 -547 545 -535
rect 745 -59 803 -47
rect 745 -535 757 -59
rect 791 -535 803 -59
rect 745 -547 803 -535
rect 1003 -59 1061 -47
rect 1003 -535 1015 -59
rect 1049 -535 1061 -59
rect 1003 -547 1061 -535
rect 1261 -59 1319 -47
rect 1261 -535 1273 -59
rect 1307 -535 1319 -59
rect 1261 -547 1319 -535
rect 1519 -59 1577 -47
rect 1519 -535 1531 -59
rect 1565 -535 1577 -59
rect 1519 -547 1577 -535
rect 1777 -59 1835 -47
rect 1777 -535 1789 -59
rect 1823 -535 1835 -59
rect 1777 -547 1835 -535
rect 2035 -59 2093 -47
rect 2035 -535 2047 -59
rect 2081 -535 2093 -59
rect 2035 -547 2093 -535
rect 2293 -59 2351 -47
rect 2293 -535 2305 -59
rect 2339 -535 2351 -59
rect 2293 -547 2351 -535
<< ndiffc >>
rect -2339 59 -2305 535
rect -2081 59 -2047 535
rect -1823 59 -1789 535
rect -1565 59 -1531 535
rect -1307 59 -1273 535
rect -1049 59 -1015 535
rect -791 59 -757 535
rect -533 59 -499 535
rect -275 59 -241 535
rect -17 59 17 535
rect 241 59 275 535
rect 499 59 533 535
rect 757 59 791 535
rect 1015 59 1049 535
rect 1273 59 1307 535
rect 1531 59 1565 535
rect 1789 59 1823 535
rect 2047 59 2081 535
rect 2305 59 2339 535
rect -2339 -535 -2305 -59
rect -2081 -535 -2047 -59
rect -1823 -535 -1789 -59
rect -1565 -535 -1531 -59
rect -1307 -535 -1273 -59
rect -1049 -535 -1015 -59
rect -791 -535 -757 -59
rect -533 -535 -499 -59
rect -275 -535 -241 -59
rect -17 -535 17 -59
rect 241 -535 275 -59
rect 499 -535 533 -59
rect 757 -535 791 -59
rect 1015 -535 1049 -59
rect 1273 -535 1307 -59
rect 1531 -535 1565 -59
rect 1789 -535 1823 -59
rect 2047 -535 2081 -59
rect 2305 -535 2339 -59
<< poly >>
rect -2293 547 -2093 573
rect -2035 547 -1835 573
rect -1777 547 -1577 573
rect -1519 547 -1319 573
rect -1261 547 -1061 573
rect -1003 547 -803 573
rect -745 547 -545 573
rect -487 547 -287 573
rect -229 547 -29 573
rect 29 547 229 573
rect 287 547 487 573
rect 545 547 745 573
rect 803 547 1003 573
rect 1061 547 1261 573
rect 1319 547 1519 573
rect 1577 547 1777 573
rect 1835 547 2035 573
rect 2093 547 2293 573
rect -2293 21 -2093 47
rect -2035 21 -1835 47
rect -1777 21 -1577 47
rect -1519 21 -1319 47
rect -1261 21 -1061 47
rect -1003 21 -803 47
rect -745 21 -545 47
rect -487 21 -287 47
rect -229 21 -29 47
rect 29 21 229 47
rect 287 21 487 47
rect 545 21 745 47
rect 803 21 1003 47
rect 1061 21 1261 47
rect 1319 21 1519 47
rect 1577 21 1777 47
rect 1835 21 2035 47
rect 2093 21 2293 47
rect -2293 -47 -2093 -21
rect -2035 -47 -1835 -21
rect -1777 -47 -1577 -21
rect -1519 -47 -1319 -21
rect -1261 -47 -1061 -21
rect -1003 -47 -803 -21
rect -745 -47 -545 -21
rect -487 -47 -287 -21
rect -229 -47 -29 -21
rect 29 -47 229 -21
rect 287 -47 487 -21
rect 545 -47 745 -21
rect 803 -47 1003 -21
rect 1061 -47 1261 -21
rect 1319 -47 1519 -21
rect 1577 -47 1777 -21
rect 1835 -47 2035 -21
rect 2093 -47 2293 -21
rect -2293 -573 -2093 -547
rect -2035 -573 -1835 -547
rect -1777 -573 -1577 -547
rect -1519 -573 -1319 -547
rect -1261 -573 -1061 -547
rect -1003 -573 -803 -547
rect -745 -573 -545 -547
rect -487 -573 -287 -547
rect -229 -573 -29 -547
rect 29 -573 229 -547
rect 287 -573 487 -547
rect 545 -573 745 -547
rect 803 -573 1003 -547
rect 1061 -573 1261 -547
rect 1319 -573 1519 -547
rect 1577 -573 1777 -547
rect 1835 -573 2035 -547
rect 2093 -573 2293 -547
<< locali >>
rect -2339 535 -2305 551
rect -2339 43 -2305 59
rect -2081 535 -2047 551
rect -2081 43 -2047 59
rect -1823 535 -1789 551
rect -1823 43 -1789 59
rect -1565 535 -1531 551
rect -1565 43 -1531 59
rect -1307 535 -1273 551
rect -1307 43 -1273 59
rect -1049 535 -1015 551
rect -1049 43 -1015 59
rect -791 535 -757 551
rect -791 43 -757 59
rect -533 535 -499 551
rect -533 43 -499 59
rect -275 535 -241 551
rect -275 43 -241 59
rect -17 535 17 551
rect -17 43 17 59
rect 241 535 275 551
rect 241 43 275 59
rect 499 535 533 551
rect 499 43 533 59
rect 757 535 791 551
rect 757 43 791 59
rect 1015 535 1049 551
rect 1015 43 1049 59
rect 1273 535 1307 551
rect 1273 43 1307 59
rect 1531 535 1565 551
rect 1531 43 1565 59
rect 1789 535 1823 551
rect 1789 43 1823 59
rect 2047 535 2081 551
rect 2047 43 2081 59
rect 2305 535 2339 551
rect 2305 43 2339 59
rect -2339 -59 -2305 -43
rect -2339 -551 -2305 -535
rect -2081 -59 -2047 -43
rect -2081 -551 -2047 -535
rect -1823 -59 -1789 -43
rect -1823 -551 -1789 -535
rect -1565 -59 -1531 -43
rect -1565 -551 -1531 -535
rect -1307 -59 -1273 -43
rect -1307 -551 -1273 -535
rect -1049 -59 -1015 -43
rect -1049 -551 -1015 -535
rect -791 -59 -757 -43
rect -791 -551 -757 -535
rect -533 -59 -499 -43
rect -533 -551 -499 -535
rect -275 -59 -241 -43
rect -275 -551 -241 -535
rect -17 -59 17 -43
rect -17 -551 17 -535
rect 241 -59 275 -43
rect 241 -551 275 -535
rect 499 -59 533 -43
rect 499 -551 533 -535
rect 757 -59 791 -43
rect 757 -551 791 -535
rect 1015 -59 1049 -43
rect 1015 -551 1049 -535
rect 1273 -59 1307 -43
rect 1273 -551 1307 -535
rect 1531 -59 1565 -43
rect 1531 -551 1565 -535
rect 1789 -59 1823 -43
rect 1789 -551 1823 -535
rect 2047 -59 2081 -43
rect 2047 -551 2081 -535
rect 2305 -59 2339 -43
rect 2305 -551 2339 -535
<< viali >>
rect -2339 59 -2305 535
rect -2081 59 -2047 535
rect -1823 59 -1789 535
rect -1565 59 -1531 535
rect -1307 59 -1273 535
rect -1049 59 -1015 535
rect -791 59 -757 535
rect -533 59 -499 535
rect -275 59 -241 535
rect -17 59 17 535
rect 241 59 275 535
rect 499 59 533 535
rect 757 59 791 535
rect 1015 59 1049 535
rect 1273 59 1307 535
rect 1531 59 1565 535
rect 1789 59 1823 535
rect 2047 59 2081 535
rect 2305 59 2339 535
rect -2339 -535 -2305 -59
rect -2081 -535 -2047 -59
rect -1823 -535 -1789 -59
rect -1565 -535 -1531 -59
rect -1307 -535 -1273 -59
rect -1049 -535 -1015 -59
rect -791 -535 -757 -59
rect -533 -535 -499 -59
rect -275 -535 -241 -59
rect -17 -535 17 -59
rect 241 -535 275 -59
rect 499 -535 533 -59
rect 757 -535 791 -59
rect 1015 -535 1049 -59
rect 1273 -535 1307 -59
rect 1531 -535 1565 -59
rect 1789 -535 1823 -59
rect 2047 -535 2081 -59
rect 2305 -535 2339 -59
<< metal1 >>
rect -2345 535 -2299 547
rect -2345 59 -2339 535
rect -2305 59 -2299 535
rect -2345 47 -2299 59
rect -2087 535 -2041 547
rect -2087 59 -2081 535
rect -2047 59 -2041 535
rect -2087 47 -2041 59
rect -1829 535 -1783 547
rect -1829 59 -1823 535
rect -1789 59 -1783 535
rect -1829 47 -1783 59
rect -1571 535 -1525 547
rect -1571 59 -1565 535
rect -1531 59 -1525 535
rect -1571 47 -1525 59
rect -1313 535 -1267 547
rect -1313 59 -1307 535
rect -1273 59 -1267 535
rect -1313 47 -1267 59
rect -1055 535 -1009 547
rect -1055 59 -1049 535
rect -1015 59 -1009 535
rect -1055 47 -1009 59
rect -797 535 -751 547
rect -797 59 -791 535
rect -757 59 -751 535
rect -797 47 -751 59
rect -539 535 -493 547
rect -539 59 -533 535
rect -499 59 -493 535
rect -539 47 -493 59
rect -281 535 -235 547
rect -281 59 -275 535
rect -241 59 -235 535
rect -281 47 -235 59
rect -23 535 23 547
rect -23 59 -17 535
rect 17 59 23 535
rect -23 47 23 59
rect 235 535 281 547
rect 235 59 241 535
rect 275 59 281 535
rect 235 47 281 59
rect 493 535 539 547
rect 493 59 499 535
rect 533 59 539 535
rect 493 47 539 59
rect 751 535 797 547
rect 751 59 757 535
rect 791 59 797 535
rect 751 47 797 59
rect 1009 535 1055 547
rect 1009 59 1015 535
rect 1049 59 1055 535
rect 1009 47 1055 59
rect 1267 535 1313 547
rect 1267 59 1273 535
rect 1307 59 1313 535
rect 1267 47 1313 59
rect 1525 535 1571 547
rect 1525 59 1531 535
rect 1565 59 1571 535
rect 1525 47 1571 59
rect 1783 535 1829 547
rect 1783 59 1789 535
rect 1823 59 1829 535
rect 1783 47 1829 59
rect 2041 535 2087 547
rect 2041 59 2047 535
rect 2081 59 2087 535
rect 2041 47 2087 59
rect 2299 535 2345 547
rect 2299 59 2305 535
rect 2339 59 2345 535
rect 2299 47 2345 59
rect -2345 -59 -2299 -47
rect -2345 -535 -2339 -59
rect -2305 -535 -2299 -59
rect -2345 -547 -2299 -535
rect -2087 -59 -2041 -47
rect -2087 -535 -2081 -59
rect -2047 -535 -2041 -59
rect -2087 -547 -2041 -535
rect -1829 -59 -1783 -47
rect -1829 -535 -1823 -59
rect -1789 -535 -1783 -59
rect -1829 -547 -1783 -535
rect -1571 -59 -1525 -47
rect -1571 -535 -1565 -59
rect -1531 -535 -1525 -59
rect -1571 -547 -1525 -535
rect -1313 -59 -1267 -47
rect -1313 -535 -1307 -59
rect -1273 -535 -1267 -59
rect -1313 -547 -1267 -535
rect -1055 -59 -1009 -47
rect -1055 -535 -1049 -59
rect -1015 -535 -1009 -59
rect -1055 -547 -1009 -535
rect -797 -59 -751 -47
rect -797 -535 -791 -59
rect -757 -535 -751 -59
rect -797 -547 -751 -535
rect -539 -59 -493 -47
rect -539 -535 -533 -59
rect -499 -535 -493 -59
rect -539 -547 -493 -535
rect -281 -59 -235 -47
rect -281 -535 -275 -59
rect -241 -535 -235 -59
rect -281 -547 -235 -535
rect -23 -59 23 -47
rect -23 -535 -17 -59
rect 17 -535 23 -59
rect -23 -547 23 -535
rect 235 -59 281 -47
rect 235 -535 241 -59
rect 275 -535 281 -59
rect 235 -547 281 -535
rect 493 -59 539 -47
rect 493 -535 499 -59
rect 533 -535 539 -59
rect 493 -547 539 -535
rect 751 -59 797 -47
rect 751 -535 757 -59
rect 791 -535 797 -59
rect 751 -547 797 -535
rect 1009 -59 1055 -47
rect 1009 -535 1015 -59
rect 1049 -535 1055 -59
rect 1009 -547 1055 -535
rect 1267 -59 1313 -47
rect 1267 -535 1273 -59
rect 1307 -535 1313 -59
rect 1267 -547 1313 -535
rect 1525 -59 1571 -47
rect 1525 -535 1531 -59
rect 1565 -535 1571 -59
rect 1525 -547 1571 -535
rect 1783 -59 1829 -47
rect 1783 -535 1789 -59
rect 1823 -535 1829 -59
rect 1783 -547 1829 -535
rect 2041 -59 2087 -47
rect 2041 -535 2047 -59
rect 2081 -535 2087 -59
rect 2041 -547 2087 -535
rect 2299 -59 2345 -47
rect 2299 -535 2305 -59
rect 2339 -535 2345 -59
rect 2299 -547 2345 -535
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 1 m 2 nf 18 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
