magic
tech sky130A
magscale 1 2
timestamp 1697926267
<< pwell >>
rect -201 -2798 201 2798
<< psubdiff >>
rect -165 2728 -69 2762
rect 69 2728 165 2762
rect -165 2666 -131 2728
rect 131 2666 165 2728
rect -165 -2728 -131 -2666
rect 131 -2728 165 -2666
rect -165 -2762 -69 -2728
rect 69 -2762 165 -2728
<< psubdiffcont >>
rect -69 2728 69 2762
rect -165 -2666 -131 2666
rect 131 -2666 165 2666
rect -69 -2762 69 -2728
<< xpolycontact >>
rect -35 2200 35 2632
rect -35 -2632 35 -2200
<< ppolyres >>
rect -35 -2200 35 2200
<< locali >>
rect -165 2728 -69 2762
rect 69 2728 165 2762
rect -165 2666 -131 2728
rect 131 2666 165 2728
rect -165 -2728 -131 -2666
rect 131 -2728 165 -2666
rect -165 -2762 -69 -2728
rect 69 -2762 165 -2728
<< viali >>
rect -19 2217 19 2614
rect -19 -2614 19 -2217
<< metal1 >>
rect -25 2614 25 2626
rect -25 2217 -19 2614
rect 19 2217 25 2614
rect -25 2205 25 2217
rect -25 -2217 25 -2205
rect -25 -2614 -19 -2217
rect 19 -2614 25 -2217
rect -25 -2626 25 -2614
<< res0p35 >>
rect -37 -2202 37 2202
<< properties >>
string FIXED_BBOX -148 -2745 148 2745
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 22.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 21.214k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
