magic
tech sky130A
magscale 1 2
timestamp 1698302399
<< nwell >>
rect 16187 -19838 23511 -19833
rect 10068 -30519 29597 -19838
<< poly >>
rect 16151 -20927 16823 -19927
rect 22875 -20927 23547 -19927
rect 16151 -21001 16823 -20985
rect 16151 -21969 16197 -21001
rect 16777 -21969 16823 -21001
rect 16151 -21985 16823 -21969
rect 22875 -21001 23547 -20985
rect 22875 -21969 22921 -21001
rect 23501 -21969 23547 -21001
rect 22875 -21985 23547 -21969
rect 16151 -22059 16823 -22043
rect 16151 -23027 16197 -22059
rect 16777 -23027 16823 -22059
rect 16151 -23043 16823 -23027
rect 22875 -22059 23547 -22043
rect 22875 -23027 22921 -22059
rect 23501 -23027 23547 -22059
rect 22875 -23043 23547 -23027
rect 16151 -23117 16823 -23101
rect 16151 -24085 16197 -23117
rect 16777 -24085 16823 -23117
rect 16151 -24101 16823 -24085
rect 22875 -23117 23547 -23101
rect 22875 -24085 22921 -23117
rect 23501 -24085 23547 -23117
rect 22875 -24101 23547 -24085
rect 16151 -24175 16823 -24159
rect 16151 -25143 16197 -24175
rect 16777 -25143 16823 -24175
rect 16151 -25159 16823 -25143
rect 22875 -24175 23547 -24159
rect 22875 -25143 22921 -24175
rect 23501 -25143 23547 -24175
rect 22875 -25159 23547 -25143
rect 16151 -25233 16823 -25217
rect 16151 -26201 16197 -25233
rect 16777 -26201 16823 -25233
rect 16151 -26217 16823 -26201
rect 22875 -25233 23547 -25217
rect 22875 -26201 22921 -25233
rect 23501 -26201 23547 -25233
rect 22875 -26217 23547 -26201
rect 16151 -26291 16823 -26275
rect 16151 -27259 16197 -26291
rect 16777 -27259 16823 -26291
rect 16151 -27275 16823 -27259
rect 22875 -26291 23547 -26275
rect 22875 -27259 22921 -26291
rect 23501 -27259 23547 -26291
rect 22875 -27275 23547 -27259
rect 16151 -27349 16823 -27333
rect 16151 -28317 16197 -27349
rect 16777 -28317 16823 -27349
rect 16151 -28333 16823 -28317
rect 22875 -27349 23547 -27333
rect 22875 -28317 22921 -27349
rect 23501 -28317 23547 -27349
rect 22875 -28333 23547 -28317
rect 16151 -28407 16823 -28391
rect 16151 -29375 16197 -28407
rect 16777 -29375 16823 -28407
rect 16151 -29391 16823 -29375
rect 22875 -28407 23547 -28391
rect 22875 -29375 22921 -28407
rect 23501 -29375 23547 -28407
rect 22875 -29391 23547 -29375
rect 16151 -30449 16823 -29449
rect 22875 -30449 23547 -29449
rect -4089 -34017 -3089 -33999
rect -4089 -34053 -4073 -34017
rect -3105 -34053 -3089 -34017
rect -4089 -34071 -3089 -34053
rect -3031 -34017 -2031 -33999
rect -3031 -34053 -3015 -34017
rect -2047 -34053 -2031 -34017
rect -3031 -34071 -2031 -34053
rect -1973 -34017 -973 -33999
rect -1973 -34053 -1957 -34017
rect -989 -34053 -973 -34017
rect -1973 -34071 -973 -34053
rect -915 -34017 85 -33999
rect -915 -34053 -899 -34017
rect 69 -34053 85 -34017
rect -915 -34071 85 -34053
rect 143 -34017 1143 -33999
rect 143 -34053 159 -34017
rect 1127 -34053 1143 -34017
rect 143 -34071 1143 -34053
rect 1201 -34017 2201 -33999
rect 1201 -34053 1217 -34017
rect 2185 -34053 2201 -34017
rect 1201 -34071 2201 -34053
rect 2259 -34017 3259 -33999
rect 2259 -34053 2275 -34017
rect 3243 -34053 3259 -34017
rect 2259 -34071 3259 -34053
rect 3317 -34017 4317 -33999
rect 3317 -34053 3333 -34017
rect 4301 -34053 4317 -34017
rect 3317 -34071 4317 -34053
rect 4375 -34017 5375 -33999
rect 4375 -34053 4391 -34017
rect 5359 -34053 5375 -34017
rect 4375 -34071 5375 -34053
rect 5433 -34017 6433 -33999
rect 5433 -34053 5449 -34017
rect 6417 -34053 6433 -34017
rect 5433 -34071 6433 -34053
<< polycont >>
rect 16197 -21969 16777 -21001
rect 22921 -21969 23501 -21001
rect 16197 -23027 16777 -22059
rect 22921 -23027 23501 -22059
rect 16197 -24085 16777 -23117
rect 22921 -24085 23501 -23117
rect 16197 -25143 16777 -24175
rect 22921 -25143 23501 -24175
rect 16197 -26201 16777 -25233
rect 22921 -26201 23501 -25233
rect 16197 -27259 16777 -26291
rect 22921 -27259 23501 -26291
rect 16197 -28317 16777 -27349
rect 22921 -28317 23501 -27349
rect 16197 -29375 16777 -28407
rect 22921 -29375 23501 -28407
rect -4073 -34053 -3105 -34017
rect -3015 -34053 -2047 -34017
rect -1957 -34053 -989 -34017
rect -899 -34053 69 -34017
rect 159 -34053 1127 -34017
rect 1217 -34053 2185 -34017
rect 2275 -34053 3243 -34017
rect 3333 -34053 4301 -34017
rect 4391 -34053 5359 -34017
rect 5449 -34053 6417 -34017
<< locali >>
rect 16181 -21001 16793 -20985
rect 16181 -21969 16197 -21001
rect 16777 -21969 16793 -21001
rect 16181 -22059 16793 -21969
rect 16181 -23027 16197 -22059
rect 16777 -23027 16793 -22059
rect 16181 -23117 16793 -23027
rect 16181 -24085 16197 -23117
rect 16777 -24085 16793 -23117
rect 16181 -24175 16793 -24085
rect 16181 -25143 16197 -24175
rect 16777 -25143 16793 -24175
rect 16181 -25233 16793 -25143
rect 16181 -26201 16197 -25233
rect 16777 -26201 16793 -25233
rect 16181 -26291 16793 -26201
rect 16181 -27259 16197 -26291
rect 16777 -27259 16793 -26291
rect 16181 -27349 16793 -27259
rect 16181 -28317 16197 -27349
rect 16777 -28317 16793 -27349
rect 16181 -28407 16793 -28317
rect 16181 -29375 16197 -28407
rect 16777 -29375 16793 -28407
rect 16181 -29391 16793 -29375
rect 22905 -21001 23517 -20985
rect 22905 -21969 22921 -21001
rect 23501 -21969 23517 -21001
rect 22905 -22059 23517 -21969
rect 22905 -23027 22921 -22059
rect 23501 -23027 23517 -22059
rect 22905 -23117 23517 -23027
rect 22905 -24085 22921 -23117
rect 23501 -24085 23517 -23117
rect 22905 -24175 23517 -24085
rect 22905 -25143 22921 -24175
rect 23501 -25143 23517 -24175
rect 22905 -25233 23517 -25143
rect 22905 -26201 22921 -25233
rect 23501 -26201 23517 -25233
rect 22905 -26291 23517 -26201
rect 22905 -27259 22921 -26291
rect 23501 -27259 23517 -26291
rect 22905 -27349 23517 -27259
rect 22905 -28317 22921 -27349
rect 23501 -28317 23517 -27349
rect 22905 -28407 23517 -28317
rect 22905 -29375 22921 -28407
rect 23501 -29375 23517 -28407
rect 22905 -29391 23517 -29375
rect -4073 -34011 -3105 -34001
rect -4073 -34017 -4063 -34011
rect -3115 -34017 -3105 -34011
rect -4073 -34059 -4063 -34053
rect -3115 -34059 -3105 -34053
rect -4073 -34069 -3105 -34059
rect -3015 -34011 -2047 -34001
rect -3015 -34017 -3005 -34011
rect -2057 -34017 -2047 -34011
rect -3015 -34059 -3005 -34053
rect -2057 -34059 -2047 -34053
rect -3015 -34069 -2047 -34059
rect -1957 -34011 -989 -34001
rect -1957 -34017 -1947 -34011
rect -999 -34017 -989 -34011
rect -1957 -34059 -1947 -34053
rect -999 -34059 -989 -34053
rect -1957 -34069 -989 -34059
rect -899 -34011 69 -34001
rect -899 -34017 -889 -34011
rect 59 -34017 69 -34011
rect -899 -34059 -889 -34053
rect 59 -34059 69 -34053
rect -899 -34069 69 -34059
rect 159 -34011 1127 -34001
rect 159 -34017 169 -34011
rect 1117 -34017 1127 -34011
rect 159 -34059 169 -34053
rect 1117 -34059 1127 -34053
rect 159 -34069 1127 -34059
rect 1217 -34011 2185 -34001
rect 1217 -34017 1227 -34011
rect 2175 -34017 2185 -34011
rect 1217 -34059 1227 -34053
rect 2175 -34059 2185 -34053
rect 1217 -34069 2185 -34059
rect 2275 -34011 3243 -34001
rect 2275 -34017 2285 -34011
rect 3233 -34017 3243 -34011
rect 2275 -34059 2285 -34053
rect 3233 -34059 3243 -34053
rect 2275 -34069 3243 -34059
rect 3333 -34011 4301 -34001
rect 3333 -34017 3343 -34011
rect 4291 -34017 4301 -34011
rect 3333 -34059 3343 -34053
rect 4291 -34059 4301 -34053
rect 3333 -34069 4301 -34059
rect 4391 -34011 5359 -34001
rect 4391 -34017 4401 -34011
rect 5349 -34017 5359 -34011
rect 4391 -34059 4401 -34053
rect 5349 -34059 5359 -34053
rect 4391 -34069 5359 -34059
rect 5449 -34011 6417 -34001
rect 5449 -34017 5459 -34011
rect 6407 -34017 6417 -34011
rect 5449 -34059 5459 -34053
rect 6407 -34059 6417 -34053
rect 5449 -34069 6417 -34059
<< viali >>
rect 16197 -21969 16777 -21001
rect 16197 -23027 16777 -22059
rect 16197 -24085 16777 -23117
rect 16197 -25143 16777 -24175
rect 16197 -26201 16777 -25233
rect 16197 -27259 16777 -26291
rect 16197 -28317 16777 -27349
rect 16197 -29375 16777 -28407
rect 22921 -21969 23501 -21001
rect 22921 -23027 23501 -22059
rect 22921 -24085 23501 -23117
rect 22921 -25143 23501 -24175
rect 22921 -26201 23501 -25233
rect 22921 -27259 23501 -26291
rect 22921 -28317 23501 -27349
rect 22921 -29375 23501 -28407
rect -4063 -34017 -3115 -34011
rect -4063 -34053 -3115 -34017
rect -4063 -34059 -3115 -34053
rect -3005 -34017 -2057 -34011
rect -3005 -34053 -2057 -34017
rect -3005 -34059 -2057 -34053
rect -1947 -34017 -999 -34011
rect -1947 -34053 -999 -34017
rect -1947 -34059 -999 -34053
rect -889 -34017 59 -34011
rect -889 -34053 59 -34017
rect -889 -34059 59 -34053
rect 169 -34017 1117 -34011
rect 169 -34053 1117 -34017
rect 169 -34059 1117 -34053
rect 1227 -34017 2175 -34011
rect 1227 -34053 2175 -34017
rect 1227 -34059 2175 -34053
rect 2285 -34017 3233 -34011
rect 2285 -34053 3233 -34017
rect 2285 -34059 3233 -34053
rect 3343 -34017 4291 -34011
rect 3343 -34053 4291 -34017
rect 3343 -34059 4291 -34053
rect 4401 -34017 5349 -34011
rect 4401 -34053 5349 -34017
rect 4401 -34059 5349 -34053
rect 5459 -34017 6407 -34011
rect 5459 -34053 6407 -34017
rect 5459 -34059 6407 -34053
<< metal1 >>
rect 16181 -21001 16793 -20985
rect 16181 -21969 16197 -21001
rect 16777 -21969 16793 -21001
rect 16181 -22059 16793 -21969
rect 16181 -23027 16197 -22059
rect 16777 -23027 16793 -22059
rect 16181 -23117 16793 -23027
rect 16181 -24085 16197 -23117
rect 16777 -24085 16793 -23117
rect 16181 -24175 16793 -24085
rect 16181 -25143 16197 -24175
rect 16777 -25143 16793 -24175
rect 16181 -25233 16793 -25143
rect 16181 -26201 16197 -25233
rect 16777 -26201 16793 -25233
rect 16181 -26291 16793 -26201
rect 16181 -27259 16197 -26291
rect 16777 -27259 16793 -26291
rect 16181 -27349 16793 -27259
rect 16181 -28317 16197 -27349
rect 16777 -28317 16793 -27349
rect 16181 -28407 16793 -28317
rect 16181 -29375 16197 -28407
rect 16777 -29375 16793 -28407
rect 16181 -29391 16793 -29375
rect 22905 -21001 23517 -20985
rect 22905 -21969 22921 -21001
rect 23501 -21969 23517 -21001
rect 22905 -22059 23517 -21969
rect 22905 -23027 22921 -22059
rect 23501 -23027 23517 -22059
rect 22905 -23117 23517 -23027
rect 22905 -24085 22921 -23117
rect 23501 -24085 23517 -23117
rect 22905 -24175 23517 -24085
rect 22905 -25143 22921 -24175
rect 23501 -25143 23517 -24175
rect 22905 -25233 23517 -25143
rect 22905 -26201 22921 -25233
rect 23501 -26201 23517 -25233
rect 22905 -26291 23517 -26201
rect 22905 -27259 22921 -26291
rect 23501 -27259 23517 -26291
rect 22905 -27349 23517 -27259
rect 22905 -28317 22921 -27349
rect 23501 -28317 23517 -27349
rect 22905 -28407 23517 -28317
rect 22905 -29375 22921 -28407
rect 23501 -29375 23517 -28407
rect 22905 -29391 23517 -29375
rect -4089 -34011 -3089 -34001
rect -4089 -34059 -4063 -34011
rect -3115 -34059 -3089 -34011
rect -4089 -34069 -3089 -34059
rect -3031 -34011 5375 -34001
rect -3031 -34059 -3005 -34011
rect -2057 -34059 -1947 -34011
rect -999 -34059 -889 -34011
rect 59 -34059 169 -34011
rect 1117 -34059 1227 -34011
rect 2175 -34059 2285 -34011
rect 3233 -34059 3343 -34011
rect 4291 -34059 4401 -34011
rect 5349 -34059 5375 -34011
rect -3031 -34069 5375 -34059
rect 5433 -34011 6433 -34001
rect 5433 -34059 5459 -34011
rect 6407 -34059 6433 -34011
rect 5433 -34069 6433 -34059
rect -4154 -37136 -4144 -36499
rect -4092 -37136 -4082 -36499
rect -2038 -37136 -2028 -36499
rect -1976 -37136 -1966 -36499
rect 78 -37136 88 -36499
rect 140 -37136 150 -36499
rect 2194 -37136 2204 -36499
rect 2256 -37136 2266 -36499
rect 4310 -37136 4320 -36499
rect 4372 -37136 4382 -36499
rect 6426 -37136 6436 -36499
rect 6488 -37136 6498 -36499
<< via1 >>
rect -4144 -37136 -4092 -36499
rect -2028 -37136 -1976 -36499
rect 88 -37136 140 -36499
rect 2204 -37136 2256 -36499
rect 4320 -37136 4372 -36499
rect 6436 -37136 6488 -36499
<< metal2 >>
rect -4141 -31581 6491 -30924
rect -4147 -33254 6485 -32597
rect -4141 -35473 6491 -34816
rect -4147 -36499 6491 -36489
rect -4147 -37136 -4144 -36499
rect -4092 -37136 -2028 -36499
rect -1976 -37136 88 -36499
rect 140 -37136 2204 -36499
rect 2256 -37136 4320 -36499
rect 4372 -37136 6436 -36499
rect 6488 -37136 6498 -36499
rect -4147 -37146 6491 -37136
use sky130_fd_pr__pfet_01v8_lvt_S6HGXS  XM1
timestamp 1697926798
transform 0 1 26573 -1 0 -25188
box -5355 -3062 5355 3062
use sky130_fd_pr__pfet_01v8_lvt_S6HGXS  XM3
timestamp 1697926798
transform 0 1 19849 -1 0 -25188
box -5355 -3062 5355 3062
use sky130_fd_pr__nfet_01v8_lvt_L9PRSH  XM11
timestamp 1698065204
transform 1 0 8237 0 1 -24815
box -558 -3088 558 3088
use sky130_fd_pr__res_high_po_0p35_N5VAUY  XR1
timestamp 1697926267
transform 1 0 -2282 0 1 -25425
box -201 -2098 201 2098
use sky130_fd_pr__res_high_po_0p35_N5VAUY  XR2
timestamp 1697926267
transform 1 0 -2684 0 1 -25425
box -201 -2098 201 2098
use sky130_fd_pr__res_high_po_0p35_N5VAUY  XR7
timestamp 1697926267
transform 1 0 -3086 0 1 -25425
box -201 -2098 201 2098
use sky130_fd_pr__res_high_po_0p35_WZDALF  XR8
timestamp 1697926267
transform 1 0 -3488 0 1 -26045
box -201 -1478 201 1478
use sky130_fd_pr__res_high_po_0p35_NBFPG6  XR9
timestamp 1697926267
transform 1 0 -3890 0 1 -25025
box -201 -2498 201 2498
use sky130_fd_pr__res_high_po_0p35_2QX5YR  XR10
timestamp 1697926267
transform 1 0 -1880 0 1 -24725
box -201 -2798 201 2798
use sky130_fd_pr__res_high_po_0p35_GF4C8W  XR11
timestamp 1697926267
transform 1 0 -1478 0 1 -24395
box -201 -3128 201 3128
use sky130_fd_pr__res_high_po_0p35_GMRRB5  XR12
timestamp 1697926267
transform 1 0 -1076 0 1 -24225
box -201 -3298 201 3298
use sky130_fd_pr__nfet_01v8_lvt_ERQKXW  sky130_fd_pr__nfet_01v8_lvt_ERQKXW_1
timestamp 1697926798
transform 1 0 1172 0 1 -37097
box -5319 -3026 5319 3026
use sky130_fd_pr__nfet_01v8_lvt_ERQKXW  sky130_fd_pr__nfet_01v8_lvt_ERQKXW_2
timestamp 1697926798
transform 1 0 1172 0 1 -30973
box -5319 -3026 5319 3026
use sky130_fd_pr__pfet_01v8_lvt_S6HGXS  sky130_fd_pr__pfet_01v8_lvt_S6HGXS_0
timestamp 1697926798
transform 0 1 13125 -1 0 -25188
box -5355 -3062 5355 3062
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1675710598
transform 0 1 3491 -1 0 -24583
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1675710598
transform 0 1 1891 -1 0 -24583
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1675710598
transform 0 1 1891 -1 0 -26183
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1675710598
transform 0 1 3491 -1 0 -26183
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1675710598
transform 0 1 5091 -1 0 -26183
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1675710598
transform 0 1 5091 -1 0 -24583
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1675710598
transform 0 1 5091 -1 0 -22983
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1675710598
transform 0 1 3491 -1 0 -22983
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1675710598
transform 0 1 1891 -1 0 -22983
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9
timestamp 1675710598
transform 0 1 3491 -1 0 -21383
box 0 0 1340 1340
use sky130_fd_sc_hd__ebufn_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1675710598
transform 0 1 85 -1 0 -24541
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  x2
timestamp 1675710598
transform 0 1 85 -1 0 -25277
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  x3
timestamp 1675710598
transform 0 1 85 -1 0 -26749
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  x4
timestamp 1675710598
transform 0 1 85 -1 0 -26013
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1675710598
transform 0 1 85 -1 0 -23168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  x6
timestamp 1675710598
transform 0 1 85 -1 0 -23628
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1675710598
transform 0 1 85 -1 0 -24088
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  x9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1675710598
transform 0 1 85 -1 0 -22892
box -38 -48 314 592
<< end >>
