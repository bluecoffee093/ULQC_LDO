* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_KPD88M w_n785_n300# a_15_n200# a_n561_n200# a_n177_n200#
+ a_111_n200# a_n129_n297# a_n513_n297# a_n609_231# a_n273_n200# a_63_n297# a_n749_n200#
+ a_687_n200# a_n321_n297# a_159_231# a_639_n297# a_n81_n200# a_399_n200# a_351_231#
+ a_495_n200# a_n33_231# a_447_n297# a_n225_231# a_591_n200# a_n657_n200# a_207_n200#
+ a_543_231# a_n369_n200# a_303_n200# a_n705_n297# a_255_n297# a_n417_231# a_n465_n200#
X0 a_n657_n200# a_n705_n297# a_n749_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X1 a_n273_n200# a_n321_n297# a_n369_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_303_n200# a_255_n297# a_207_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_591_n200# a_543_231# a_495_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_n177_n200# a_n225_231# a_n273_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X5 a_207_n200# a_159_231# a_111_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_495_n200# a_447_n297# a_399_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_n561_n200# a_n609_231# a_n657_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X8 a_111_n200# a_63_n297# a_15_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X9 a_399_n200# a_351_231# a_303_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 a_n465_n200# a_n513_n297# a_n561_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X11 a_687_n200# a_639_n297# a_591_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X12 a_n81_n200# a_n129_n297# a_n177_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X13 a_15_n200# a_n33_231# a_n81_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 a_n369_n200# a_n417_231# a_n465_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt power_transistor VDD EA_OUT BIAS_CURR OUT
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT BIAS_CURR VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT BIAS_CURR VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_A3UXRA a_3423_n1000# a_4623_1130# a_1743_1130#
+ a_3135_n1000# a_1503_n3218# a_n3297_1218# a_n4641_1218# a_1215_n3218# a_n1761_1218#
+ a_207_1130# a_n4161_n3218# a_n33_n3218# a_n3921_n1088# a_1119_1218# a_n2289_1022#
+ a_n3345_n1088# a_n3633_1022# a_4239_1130# a_1359_1130# a_3231_n1000# a_n4257_1218#
+ a_2703_1130# a_1311_n3218# a_n1377_1218# a_1023_n3218# a_n2721_1218# a_n465_3240#
+ a_n3249_1022# a_n1713_1022# a_n3153_n1088# a_2319_1130# a_n3969_n1000# a_n2337_1218#
+ a_n1329_1022# a_n4209_1022# a_n3777_n1000# a_n3489_n1000# a_n1857_n3218# a_n1569_n3218#
+ a_n609_n3218# a_n3873_n1000# a_n3585_n1000# a_n1953_n3218# a_n3297_n1000# a_n1665_n3218#
+ a_n1377_n3218# a_n1089_n3218# a_n705_n3218# a_n129_n3218# a_n417_n3218# a_n513_1218#
+ a_n3681_n1000# a_n3393_n1000# a_n1761_n3218# a_n1185_n3218# a_n1473_n3218# a_n753_1130#
+ a_3471_1022# a_n801_n3218# a_n513_n3218# a_4095_1218# a_n129_1218# a_n225_n3218#
+ a_n369_1130# a_3087_1022# a_4431_1022# a_n1281_n3218# a_1551_1022# a_n2385_3240#
+ a_n321_n3218# a_2175_1218# a_4047_1022# a_2799_n1196# a_1167_1022# a_2511_1022#
+ a_n3345_3240# a_3135_1218# a_2127_1022# a_n3393_1218# a_n4305_3240# a_n1425_3240#
+ a_1215_1218# a_2991_n1196# a_63_1218# a_n4353_1218# a_n1473_1218# a_n3729_n1196#
+ a_n4593_1130# a_n1089_1218# a_n2433_1218# a_15_1022# a_n3537_n1196# a_n2673_1130#
+ a_2895_n3306# a_4767_n3218# a_4479_n3218# a_n2049_1218# a_n3921_n1196# a_n4829_1218#
+ a_n2289_1130# a_n3345_n1196# a_n3633_1130# a_n561_1022# a_4575_n3218# a_4287_n3218#
+ a_n3009_1218# a_3183_3240# a_3759_n1088# a_n3249_1130# a_n177_1022# a_n3153_n1196#
+ a_111_3240# a_n1713_1130# a_4671_n3218# a_4383_n3218# a_4095_n3218# a_879_3240#
+ a_n3825_n3306# a_927_n3218# a_4143_3240# a_3567_n1088# a_n3249_n3306# a_639_n3218#
+ a_1263_3240# a_n4209_1130# a_n1329_1130# a_4191_n3218# a_4191_1218# a_n225_1218#
+ a_3951_n1088# a_n3633_n3306# a_735_n3218# a_2223_3240# a_n3057_n3306# a_447_n3218#
+ a_3375_n1088# a_159_n3218# a_2271_1218# a_n3441_n3306# a_831_n3218# a_543_n3218#
+ a_255_n3218# a_3183_n1088# a_3999_n1000# a_3231_1218# a_351_n3218# a_3471_1130#
+ a_3999_1218# a_n4305_n1088# a_927_1218# a_1887_n3218# a_1599_n3218# a_1311_1218#
+ a_n2481_1022# a_3087_1130# a_4431_1130# a_1551_1130# a_n4113_n1088# a_1983_n3218#
+ a_1695_n3218# a_n2097_1022# a_n3441_1022# a_63_n1000# a_4047_1130# a_2511_1130#
+ a_1167_1130# a_n1185_1218# a_n4065_1218# a_n273_3240# a_1791_n3218# a_n3057_1022#
+ a_n4737_n1000# a_n4401_1022# a_n1521_1022# a_n4449_n1000# a_n2817_n3218# a_2127_1130#
+ a_n2529_n3218# a_n2145_1218# a_n4017_1022# a_n1137_1022# a_n4545_n1000# a_n4257_n1000#
+ a_n2913_n3218# a_n2337_n3218# a_n2625_n3218# a_n3105_1218# a_n2049_n3218# a_n1809_n1088#
+ a_n4641_n1000# a_1407_n1000# a_n4353_n1000# a_1119_n1000# a_n2721_n3218# a_n4065_n1000#
+ a_n2433_n3218# a_n2145_n3218# a_15_1130# a_n1617_n1088# a_1503_n1000# a_1215_n1000#
+ a_n4161_n1000# a_n2241_n3218# a_n33_n1000# a_n321_1218# a_n897_n3218# a_n1425_n1088#
+ a_n561_1130# a_1023_n1000# a_1311_n1000# a_3759_n1196# a_975_1022# a_n993_n3218#
+ a_n177_1130# a_n1233_n1088# a_n2193_3240# a_3567_n1196# a_n1041_n1088# a_n3153_3240#
+ a_n1857_n1000# a_3951_n1196# a_n1569_n1000# a_3375_n1196# a_n609_n1000# a_n4113_3240#
+ a_639_1218# a_n1233_3240# a_n1953_n1000# a_n1665_n1000# a_n1377_n1000# a_1023_1218#
+ a_n1089_n1000# a_3183_n1196# a_n705_n1000# a_n417_n1000# a_n1281_1218# a_n4161_1218#
+ a_n129_n1000# a_3855_n3306# a_n1761_n1000# a_3279_n3306# a_n1473_n1000# a_n1185_n1000#
+ a_15_n3306# a_n801_n1000# a_n4305_n1196# a_n513_n1000# a_n225_n1000# a_n2241_1218#
+ a_3663_n3306# a_n2481_1130# a_n1281_n1000# a_3087_n3306# a_4719_n1088# a_n321_n1000#
+ a_n4113_n1196# a_n3201_1218# a_3471_n3306# a_n2097_1130# a_n3969_1218# a_n3441_1130#
+ a_4527_n1088# a_n4209_n3306# a_n3057_1130# a_n4401_1130# a_n1521_1130# a_4335_n1088#
+ a_n4017_n3306# a_687_3240# a_1071_3240# a_n4017_1130# a_n1137_1130# a_n4401_n3306#
+ a_4143_n1088# a_n1809_n1196# a_2031_3240# a_2799_3240# a_n1617_n1196# a_4479_n1000#
+ a_4767_n1000# a_2847_n3218# a_2559_n3218# a_3759_3240# a_n1425_n1196# a_n4689_n1088#
+ a_303_n1088# a_4575_n1000# a_2943_n3218# a_4719_3240# a_4287_n1000# a_2655_n3218#
+ a_1839_3240# a_2367_n3218# a_2079_n3218# a_735_1218# a_1839_n1088# a_n33_1218# a_n1233_n1196#
+ a_n4497_n1088# a_975_1130# a_111_n1088# a_4671_n1000# a_4767_1218# a_4383_n1000#
+ a_2751_n3218# a_1887_1218# a_927_n1000# a_4095_n1000# a_2463_n3218# a_639_n1000#
+ a_n1905_n3306# a_2175_n3218# a_n1329_n3306# a_1647_n1088# a_n1041_n1196# a_4191_n1000#
+ a_2847_1218# a_2271_n3218# a_447_n1000# a_735_n1000# a_n1713_n3306# a_159_n1000#
+ a_1455_n1088# a_n1137_n3306# a_n3009_n3218# a_3807_1218# a_831_n1000# a_543_n1000#
+ a_255_n1000# a_n1521_n3306# a_1263_n1088# a_n3105_n3218# a_n81_n1088# a_351_n1000#
+ a_1071_n1088# a_n3201_n3218# a_n81_3240# a_1599_n1000# a_1887_n1000# a_4719_n1196#
+ a_n849_3240# a_1983_n1000# a_1695_n1000# a_n849_n1088# a_n897_1218# a_4527_n1196#
+ a_1791_n1000# a_n2001_n1088# a_n657_n1088# a_783_1022# a_n2817_n1000# a_n2529_n1000#
+ a_4335_n1196# a_399_1022# a_n2913_n1000# a_n465_n1088# a_n2625_n1000# a_n2337_n1000#
+ a_n2049_n1000# a_4143_n1196# a_831_1218# a_2895_1022# a_n273_n1088# a_n2721_n1000#
+ a_n2433_n1000# a_4239_n3306# a_1983_1218# a_n2145_n1000# a_n1041_3240# a_447_1218#
+ a_3855_1022# a_n4689_3240# a_4623_n3306# a_4479_1218# a_1599_1218# a_4047_n3306#
+ a_2943_1218# a_n2241_n1000# a_n2001_3240# a_n4689_n1196# a_n897_n1000# a_303_n1196#
+ a_1935_1022# a_n2769_3240# a_4431_n3306# a_3903_1218# a_2559_1218# a_1839_n1196#
+ a_n993_n1000# a_n4497_n1196# a_n3729_3240# a_111_n1196# a_3519_1218# a_1647_n1196#
+ a_207_n3306# a_n3777_1218# a_n1809_3240# a_1455_n1196# a_n4829_n3218# a_n4737_1218#
+ a_n1857_1218# a_495_3240# a_n4785_n3306# a_1263_n1196# a_n2817_1218# a_n993_1218#
+ a_2991_3240# a_n81_n1196# a_1935_n3306# a_3807_n3218# a_n4593_n3306# a_1359_n3306#
+ a_3519_n3218# a_1071_n1196# a_879_n1088# a_3951_3240# a_1743_n3306# a_n945_1022#
+ a_3903_n3218# a_3615_n3218# a_1167_n3306# a_3327_n3218# a_3039_n3218# a_3567_3240#
+ a_687_n1088# a_n849_n1196# a_1551_n3306# a_3711_n3218# a_3423_n3218# a_3135_n3218#
+ a_4527_3240# a_2607_n1088# a_1647_3240# a_495_n1088# a_n2001_n1196# a_543_1218#
+ a_n657_n1196# a_783_1130# a_3231_n3218# a_4575_1218# a_1695_1218# a_n609_1218# a_2415_n1088#
+ a_2607_3240# a_159_1218# a_399_1130# a_n465_n1196# a_n3969_n3218# a_2655_1218# a_2223_n1088#
+ a_2895_1130# a_n273_n1196# a_3615_1218# a_n3489_n3218# a_n3777_n3218# a_n4785_1022#
+ a_2031_n1088# a_n945_n3306# a_3855_1130# a_2847_n1000# a_n369_n3306# a_n3873_1218#
+ a_2559_n1000# a_n3873_n3218# a_n2865_1022# a_n3585_n3218# a_n3297_n3218# a_n2769_n1088#
+ a_1935_1130# a_n753_n3306# a_n3489_1218# a_2655_n1000# a_2943_n1000# a_n177_n3306#
+ a_n1953_1218# a_2367_n1000# a_2079_n1000# a_n3681_n3218# a_n3393_n3218# a_n3825_1022#
+ a_n4449_1218# a_n2577_n1088# a_n561_n3306# a_n1569_1218# a_n2913_1218# a_n657_3240#
+ a_2751_n1000# a_2175_n1000# a_2463_n1000# a_n1905_1022# a_n2961_n1088# a_n2529_1218#
+ a_n2385_n1088# a_2271_n1000# a_n3009_n1000# a_591_1022# a_n2193_n1088# a_n3105_n1000#
+ a_n3201_n1000# a_879_n1196# a_4671_1218# a_1791_1218# a_n705_1218# a_255_1218# a_n945_1130#
+ a_3663_1022# a_n4497_3240# a_n2961_3240# a_4287_1218# a_687_n1196# a_2751_1218#
+ a_3279_1022# a_4623_1022# a_1743_1022# a_n2577_3240# a_n3921_3240# a_207_1022# a_2607_n1196#
+ a_2367_1218# a_495_n1196# a_3711_1218# a_4239_1022# a_1359_1022# a_2703_1022# a_n3537_3240#
+ a_2415_n1196# a_3327_1218# a_2319_1022# a_n3585_1218# a_975_n3306# a_n1617_3240#
+ a_399_n3306# a_2223_n1196# a_1407_1218# a_n4545_1218# a_n1665_1218# a_783_n3306#
+ a_2319_n3306# a_n4785_1130# a_2031_n1196# a_2703_n3306# a_n2625_1218# a_591_n3306#
+ a_2127_n3306# a_n2865_1130# a_n2769_n1196# a_3999_n3218# a_2511_n3306# a_n3825_1130#
+ a_n753_1022# a_n2577_n1196# a_3375_3240# a_n369_1022# a_303_3240# a_n1905_1130#
+ a_n2961_n1196# a_n2385_n1196# a_n801_1218# a_4335_3240# a_1455_3240# a_351_1218#
+ a_n4829_n1000# a_2799_n1088# a_63_n3218# a_591_1130# a_n2193_n1196# a_4383_1218#
+ a_n417_1218# a_2415_3240# a_n2865_n3306# a_n4737_n3218# a_n2289_n3306# a_n4449_n3218#
+ a_2463_1218# a_3807_n1000# a_3519_n1000# a_n2673_n3306# a_2991_n1088# a_n4545_n3218#
+ a_n2097_n3306# a_n4257_n3218# a_2079_1218# a_n3729_n1088# a_n4593_1022# a_3423_1218#
+ a_3903_n1000# a_3327_n1000# a_3615_n1000# a_3663_1130# a_3039_n1000# a_1407_n3218#
+ VSUBS a_n2481_n3306# a_n4641_n3218# a_1119_n3218# a_n3681_1218# a_n4065_n3218# a_n4353_n3218#
+ a_3039_1218# a_n3537_n1088# a_1503_1218# a_n2673_1022# a_3711_n1000# a_3279_1130#
X0 a_n321_1218# a_n369_1130# a_n417_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X1 a_2463_n1000# a_2415_n1088# a_2367_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X2 a_n2529_1218# a_n2577_3240# a_n2625_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X3 a_3135_n3218# a_3087_n3306# a_3039_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X4 a_1119_n3218# a_1071_n1196# a_1023_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X5 a_3519_1218# a_3471_1130# a_3423_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X6 a_3135_n1000# a_3087_1022# a_3039_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X7 a_n4641_1218# a_n4689_3240# a_n4737_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X8 a_1503_1218# a_1455_3240# a_1407_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X9 a_n4257_n1000# a_n4305_n1088# a_n4353_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X10 a_1119_n1000# a_1071_n1088# a_1023_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X11 a_n129_n3218# a_n177_n3306# a_n225_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X12 a_543_1218# a_495_3240# a_447_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X13 a_159_n1000# a_111_n1088# a_63_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X14 a_1599_n3218# a_1551_n3306# a_1503_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X15 a_447_n3218# a_399_n3306# a_351_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X16 a_n1185_1218# a_n1233_3240# a_n1281_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X17 a_n2241_n1000# a_n2289_1022# a_n2337_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X18 a_2175_1218# a_2127_1130# a_2079_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X19 a_n3777_n1000# a_n3825_1022# a_n3873_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X20 a_2175_n3218# a_2127_n3306# a_2079_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X21 a_n609_n3218# a_n657_n1196# a_n705_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X22 a_4767_n1000# a_4719_n1088# a_4671_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.1e+12p pd=2.062e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X23 a_n1089_n3218# a_n1137_n3306# a_n1185_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X24 a_n2817_1218# a_n2865_1130# a_n2913_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X25 a_n225_n1000# a_n273_n1088# a_n321_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X26 a_2751_n1000# a_2703_1022# a_2655_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X27 a_4287_n3218# a_4239_n3306# a_4191_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X28 a_3807_1218# a_3759_3240# a_3711_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X29 a_2655_n3218# a_2607_n1196# a_2559_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X30 a_n3489_1218# a_n3537_3240# a_n3585_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X31 a_1791_1218# a_1743_1130# a_1695_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X32 a_1215_n3218# a_1167_n3306# a_1119_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X33 a_831_1218# a_783_1130# a_735_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X34 a_4479_1218# a_4431_1130# a_4383_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X35 a_n4545_n1000# a_n4593_1022# a_n4641_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X36 a_1407_n1000# a_1359_1022# a_1311_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X37 a_4767_n3218# a_4719_n1196# a_4671_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.1e+12p pd=2.062e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X38 a_3231_n3218# a_3183_n1196# a_3135_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X39 a_n1473_1218# a_n1521_1130# a_n1569_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X40 a_447_n1000# a_399_1022# a_351_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X41 a_2463_1218# a_2415_3240# a_2367_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X42 a_n1089_n1000# a_n1137_1022# a_n1185_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X43 a_3327_n3218# a_3279_n3306# a_3231_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X44 a_2079_n1000# a_2031_n1088# a_1983_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X45 a_1695_n3218# a_1647_n1196# a_1599_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X46 a_n225_n3218# a_n273_n1196# a_n321_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X47 a_543_n3218# a_495_n1196# a_447_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X48 a_3135_1218# a_3087_1130# a_3039_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X49 a_n3201_n1000# a_n3249_1022# a_n3297_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X50 a_n4257_1218# a_n4305_3240# a_n4353_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X51 a_1119_1218# a_1071_3240# a_1023_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X52 a_4191_n1000# a_4143_n1088# a_4095_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X53 a_3807_n3218# a_3759_n1196# a_3711_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X54 a_2271_n3218# a_2223_n1196# a_2175_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X55 a_159_1218# a_111_3240# a_63_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X56 a_n513_n1000# a_n561_1022# a_n609_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X57 a_n705_n3218# a_n753_n3306# a_n801_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X58 a_n2241_1218# a_n2289_1130# a_n2337_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X59 a_n1185_n3218# a_n1233_n1196# a_n1281_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X60 a_63_n1000# a_15_1022# a_n33_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X61 a_4383_n3218# a_4335_n1196# a_4287_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X62 a_n3777_1218# a_n3825_1130# a_n3873_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X63 a_1695_n1000# a_1647_n1088# a_1599_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X64 a_2751_n3218# a_2703_n3306# a_2655_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X65 a_4767_1218# a_4719_3240# a_4671_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.1e+12p pd=2.062e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X66 a_735_n1000# a_687_n1088# a_639_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X67 a_n3297_n3218# a_n3345_n1196# a_n3393_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X68 a_n1377_n1000# a_n1425_n1088# a_n1473_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X69 a_n225_1218# a_n273_3240# a_n321_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X70 a_2751_1218# a_2703_1130# a_2655_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X71 a_2367_n1000# a_2319_1022# a_2271_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X72 a_1311_n3218# a_1263_n1196# a_1215_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X73 a_n3777_n3218# a_n3825_n3306# a_n3873_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X74 a_3039_n1000# a_2991_n1088# a_2943_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X75 a_3423_n3218# a_3375_n1196# a_3327_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X76 a_n321_n3218# a_n369_n3306# a_n417_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X77 a_n4545_1218# a_n4593_1130# a_n4641_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X78 a_1407_1218# a_1359_1130# a_1311_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X79 a_n801_n1000# a_n849_n1088# a_n897_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X80 a_1791_n3218# a_1743_n3306# a_1695_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X81 a_n2337_n3218# a_n2385_n1196# a_n2433_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X82 a_447_1218# a_399_1130# a_351_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X83 a_n1089_1218# a_n1137_1130# a_n1185_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X84 a_n2145_n1000# a_n2193_n1088# a_n2241_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X85 a_3999_n1000# a_3951_n1088# a_3903_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X86 a_2079_1218# a_2031_3240# a_1983_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X87 a_n4449_n3218# a_n4497_n1196# a_n4545_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X88 a_3903_n3218# a_3855_n3306# a_3807_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X89 a_n801_n3218# a_n849_n1196# a_n897_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X90 a_1983_n1000# a_1935_1022# a_1887_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X91 a_n1281_n3218# a_n1329_n3306# a_n1377_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X92 a_n2817_n3218# a_n2865_n3306# a_n2913_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X93 a_n3201_1218# a_n3249_1130# a_n3297_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X94 a_4191_1218# a_4143_3240# a_4095_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X95 a_n513_1218# a_n561_1130# a_n609_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X96 a_n129_n1000# a_n177_1022# a_n225_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X97 a_2655_n1000# a_2607_n1088# a_2559_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X98 a_n3393_n3218# a_n3441_n3306# a_n3489_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X99 a_63_1218# a_15_1130# a_n33_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X100 a_1695_1218# a_1647_3240# a_1599_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X101 a_n1761_n1000# a_n1809_n1088# a_n1857_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X102 a_735_1218# a_687_3240# a_639_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X103 a_n4449_n1000# a_n4497_n1088# a_n4545_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X104 a_n1857_n3218# a_n1905_n3306# a_n1953_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X105 a_n3873_n3218# a_n3921_n1196# a_n3969_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X106 a_n1377_1218# a_n1425_3240# a_n1473_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X107 a_2367_1218# a_2319_1130# a_2271_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X108 a_n2433_n1000# a_n2481_1022# a_n2529_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X109 a_n4065_n3218# a_n4113_n1196# a_n4161_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X110 a_3423_n1000# a_3375_n1088# a_3327_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X111 a_n2433_n3218# a_n2481_n3306# a_n2529_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X112 a_n3969_n3218# a_n4017_n3306# a_n4065_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X113 a_3039_1218# a_2991_3240# a_2943_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X114 a_n3105_n1000# a_n3153_n1088# a_n3201_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X115 a_n801_1218# a_n849_3240# a_n897_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X116 a_2943_n1000# a_2895_1022# a_2847_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X117 a_4095_n1000# a_4047_1022# a_3999_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X118 a_n4545_n3218# a_n4593_n3306# a_n4641_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X119 a_n417_n1000# a_n465_n1088# a_n513_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X120 a_n2913_n3218# a_n2961_n1196# a_n3009_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X121 a_n2145_1218# a_n2193_3240# a_n2241_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X122 a_3999_1218# a_3951_3240# a_3903_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X123 a_1983_1218# a_1935_1130# a_1887_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X124 a_n4737_n1000# a_n4785_1022# a_n4829_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.1e+12p ps=2.062e+07u w=1e+07u l=150000u
X125 a_1599_n1000# a_1551_1022# a_1503_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X126 a_n2721_n1000# a_n2769_n1088# a_n2817_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X127 a_639_n1000# a_591_1022# a_543_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X128 a_n129_1218# a_n177_1130# a_n225_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X129 a_2655_1218# a_2607_3240# a_2559_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X130 a_3711_n1000# a_3663_1022# a_3615_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X131 a_n1953_n3218# a_n2001_n1196# a_n2049_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X132 a_n3393_n1000# a_n3441_1022# a_n3489_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X133 a_n4161_n3218# a_n4209_n3306# a_n4257_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X134 a_n1761_1218# a_n1809_3240# a_n1857_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X135 a_4383_n1000# a_4335_n1088# a_4287_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X136 a_n4449_1218# a_n4497_3240# a_n4545_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X137 a_n705_n1000# a_n753_1022# a_n801_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X138 a_159_n3218# a_111_n1196# a_63_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X139 a_n2433_1218# a_n2481_1130# a_n2529_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X140 a_n4641_n3218# a_n4689_n1196# a_n4737_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X141 a_63_n3218# a_15_n3306# a_n33_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X142 a_3423_1218# a_3375_3240# a_3327_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X143 a_n2049_n1000# a_n2097_1022# a_n2145_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X144 a_1887_n1000# a_1839_n1088# a_1791_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X145 a_639_n3218# a_591_n3306# a_543_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X146 a_n3105_1218# a_n3153_3240# a_n3201_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X147 a_2943_1218# a_2895_1130# a_2847_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X148 a_4095_1218# a_4047_1130# a_3999_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X149 a_n4161_n1000# a_n4209_1022# a_n4257_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X150 a_n417_1218# a_n465_3240# a_n513_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X151 a_2559_n1000# a_2511_1022# a_2463_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X152 a_2367_n3218# a_2319_n3306# a_2271_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X153 a_n3681_n1000# a_n3729_n1088# a_n3777_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X154 a_1023_n1000# a_975_1022# a_927_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X155 a_n4737_1218# a_n4785_1130# a_n4829_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.1e+12p ps=2.062e+07u w=1e+07u l=150000u
X156 a_1599_1218# a_1551_1130# a_1503_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X157 a_n1665_n1000# a_n1713_1022# a_n1761_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X158 a_4671_n1000# a_4623_1022# a_4575_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X159 a_4479_n3218# a_4431_n3306# a_4383_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X160 a_2847_n3218# a_2799_n1196# a_2751_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X161 a_n2721_1218# a_n2769_3240# a_n2817_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X162 a_639_1218# a_591_1130# a_543_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X163 a_3711_1218# a_3663_1130# a_3615_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X164 a_n2337_n1000# a_n2385_n1088# a_n2433_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X165 a_3327_n1000# a_3279_1022# a_3231_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X166 a_1407_n3218# a_1359_n3306# a_1311_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X167 a_255_n3218# a_207_n3306# a_159_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X168 a_n3393_1218# a_n3441_1130# a_n3489_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X169 a_4383_1218# a_4335_3240# a_4287_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X170 a_n3009_n1000# a_n3057_1022# a_n3105_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X171 a_1311_n1000# a_1263_n1088# a_1215_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X172 a_n705_1218# a_n753_1130# a_n801_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X173 a_351_n1000# a_303_n1088# a_255_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X174 a_2847_n1000# a_2799_n1088# a_2751_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X175 a_3519_n3218# a_3471_n3306# a_3423_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X176 a_n417_n3218# a_n465_n1196# a_n513_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X177 a_n3969_n1000# a_n4017_1022# a_n4065_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X178 a_n993_n1000# a_n1041_n1088# a_n1089_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X179 a_n33_n1000# a_n81_n1088# a_n129_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X180 a_1887_n3218# a_1839_n1196# a_1791_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X181 a_735_n3218# a_687_n1196# a_639_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X182 a_n2049_1218# a_n2097_1130# a_n2145_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X183 a_n1953_n1000# a_n2001_n1088# a_n2049_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X184 a_4095_n3218# a_4047_n3306# a_3999_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X185 a_1887_1218# a_1839_3240# a_1791_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X186 a_3999_n3218# a_3951_n1196# a_3903_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X187 a_2463_n3218# a_2415_n1196# a_2367_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X188 a_n897_n3218# a_n945_n3306# a_n993_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X189 a_n3009_n3218# a_n3057_n3306# a_n3105_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X190 a_n1377_n3218# a_n1425_n1196# a_n1473_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X191 a_n4161_1218# a_n4209_1130# a_n4257_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X192 a_2559_1218# a_2511_1130# a_2463_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X193 a_n2625_n1000# a_n2673_1022# a_n2721_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X194 a_3615_n1000# a_3567_n1088# a_3519_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X195 a_4575_n3218# a_4527_n1196# a_4479_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X196 a_2943_n3218# a_2895_n3306# a_2847_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X197 a_n3489_n3218# a_n3537_n1196# a_n3585_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X198 a_n3681_1218# a_n3729_3240# a_n3777_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X199 a_1023_1218# a_975_1130# a_927_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X200 a_n1665_1218# a_n1713_1130# a_n1761_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X201 a_4671_1218# a_4623_1130# a_4575_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X202 a_n3297_n1000# a_n3345_n1088# a_n3393_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X203 a_1503_n3218# a_1455_n1196# a_1407_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X204 a_n609_n1000# a_n657_n1088# a_n705_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X205 a_4287_n1000# a_4239_1022# a_4191_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X206 a_351_n3218# a_303_n1196# a_255_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X207 a_n2049_n3218# a_n2097_n3306# a_n2145_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X208 a_n1281_n1000# a_n1329_1022# a_n1377_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X209 a_n2337_1218# a_n2385_3240# a_n2433_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X210 a_2271_n1000# a_2223_n1088# a_2175_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X211 a_3615_n3218# a_3567_n1196# a_3519_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X212 a_3327_1218# a_3279_1130# a_3231_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X213 a_1983_n3218# a_1935_n3306# a_1887_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X214 a_n513_n3218# a_n561_n3306# a_n609_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X215 a_831_n3218# a_783_n3306# a_735_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X216 a_n993_n3218# a_n1041_n1196# a_n1089_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X217 a_n2529_n3218# a_n2577_n1196# a_n2625_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X218 a_n3009_1218# a_n3057_1130# a_n3105_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X219 a_1311_1218# a_1263_3240# a_1215_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X220 a_4191_n3218# a_4143_n1196# a_4095_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X221 a_351_1218# a_303_3240# a_255_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X222 a_2847_1218# a_2799_3240# a_2751_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X223 a_n4065_n1000# a_n4113_n1088# a_n4161_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X224 a_n2913_n1000# a_n2961_n1088# a_n3009_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X225 a_927_n3218# a_879_n1196# a_831_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X226 a_n3969_1218# a_n4017_1130# a_n4065_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X227 a_n993_1218# a_n1041_3240# a_n1089_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X228 a_n33_1218# a_n81_3240# a_n129_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X229 a_3903_n1000# a_3855_1022# a_3807_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X230 a_n3105_n3218# a_n3153_n1196# a_n3201_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X231 a_n1473_n3218# a_n1521_n3306# a_n1569_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X232 a_n1953_1218# a_n2001_3240# a_n2049_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X233 a_n3585_n1000# a_n3633_1022# a_n3681_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X234 a_927_n1000# a_879_n1088# a_831_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X235 a_4671_n3218# a_4623_n3306# a_4575_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X236 a_n1569_n1000# a_n1617_n1088# a_n1665_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.066e+07u as=0p ps=0u w=1e+07u l=150000u
X237 a_4575_n1000# a_4527_n1088# a_4479_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X238 a_n1569_n3218# a_n1617_n1196# a_n1665_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X239 a_n897_n1000# a_n945_1022# a_n993_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X240 a_n3585_n3218# a_n3633_n3306# a_n3681_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X241 a_n2625_1218# a_n2673_1130# a_n2721_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X242 a_3615_1218# a_3567_3240# a_3519_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X243 a_n2145_n3218# a_n2193_n1196# a_n2241_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X244 a_3231_n1000# a_3183_n1088# a_3135_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X245 a_n3297_1218# a_n3345_3240# a_n3393_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X246 a_n4353_n1000# a_n4401_1022# a_n4449_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X247 a_1215_n1000# a_1167_1022# a_1119_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X248 a_3711_n3218# a_3663_n3306# a_3615_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X249 a_n4257_n3218# a_n4305_n1196# a_n4353_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X250 a_n609_1218# a_n657_3240# a_n705_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X251 a_4287_1218# a_4239_1130# a_4191_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X252 a_255_n1000# a_207_1022# a_159_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X253 a_n2625_n3218# a_n2673_n3306# a_n2721_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X254 a_n1281_1218# a_n1329_1130# a_n1377_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X255 a_2271_1218# a_2223_3240# a_2175_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X256 a_1023_n3218# a_975_n3306# a_927_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X257 a_n3873_n1000# a_n3921_n1088# a_n3969_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X258 a_n4737_n3218# a_n4785_n3306# a_n4829_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.1e+12p ps=2.062e+07u w=1e+07u l=150000u
X259 a_n3201_n3218# a_n3249_n3306# a_n3297_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X260 a_n1857_n1000# a_n1905_1022# a_n1953_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X261 a_n4065_1218# a_n4113_3240# a_n4161_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X262 a_n2913_1218# a_n2961_3240# a_n3009_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X263 a_n321_n1000# a_n369_1022# a_n417_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X264 a_3903_1218# a_3855_1130# a_3807_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X265 a_n2529_n1000# a_n2577_n1088# a_n2625_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X266 a_n1665_n3218# a_n1713_n3306# a_n1761_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+12p ps=2.066e+07u w=1e+07u l=150000u
X267 a_n3681_n3218# a_n3729_n1196# a_n3777_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X268 a_3519_n1000# a_3471_1022# a_3423_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X269 a_n3585_1218# a_n3633_1130# a_n3681_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X270 a_927_1218# a_879_3240# a_831_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X271 a_n1569_1218# a_n1617_3240# a_n1665_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X272 a_4575_1218# a_4527_3240# a_4479_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X273 a_n4641_n1000# a_n4689_n1088# a_n4737_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X274 a_1503_n1000# a_1455_n1088# a_1407_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X275 a_n2241_n3218# a_n2289_n3306# a_n2337_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X276 a_n897_1218# a_n945_1130# a_n993_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X277 a_543_n1000# a_495_n1088# a_447_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X278 a_3039_n3218# a_2991_n1196# a_2943_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X279 a_n1185_n1000# a_n1233_n1088# a_n1281_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X280 a_2175_n1000# a_2127_1022# a_2079_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X281 a_n4353_n3218# a_n4401_n3306# a_n4449_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X282 a_n2721_n3218# a_n2769_n1196# a_n2817_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X283 a_3231_1218# a_3183_3240# a_3135_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X284 a_n4353_1218# a_n4401_1130# a_n4449_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X285 a_1215_1218# a_1167_1130# a_1119_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X286 a_255_1218# a_207_1130# a_159_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X287 a_n2817_n1000# a_n2865_1022# a_n2913_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X288 a_2079_n3218# a_2031_n1196# a_1983_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X289 a_3807_n1000# a_3759_n1088# a_3711_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X290 a_n33_n3218# a_n81_n1196# a_n129_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X291 a_n3873_1218# a_n3921_3240# a_n3969_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X292 a_n3489_n1000# a_n3537_n1088# a_n3585_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X293 a_1791_n1000# a_1743_1022# a_1695_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X294 a_n1761_n3218# a_n1809_n1196# a_n1857_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X295 a_n1857_1218# a_n1905_1130# a_n1953_1218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X296 a_831_n1000# a_783_1022# a_735_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X297 a_4479_n1000# a_4431_1022# a_4383_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X298 a_2559_n3218# a_2511_n3306# a_2463_n3218# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X299 a_n1473_n1000# a_n1521_1022# a_n1569_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_477Z4B a_n682_n597# a_n501_n500# a_n855_n500# a_561_n500#
+ a_n383_n500# a_n210_n597# a_n564_n597# a_n737_n500# a_797_n500# a_443_n500# a_380_n597#
+ a_n92_n597# a_n265_n500# a_n446_n597# a_734_n597# a_n619_n500# a_325_n500# a_679_n500#
+ a_n147_n500# a_262_n597# a_n328_n597# a_616_n597# w_n993_n719# a_207_n500# a_144_n597#
+ a_498_n597# a_n29_n500# a_89_n500# a_n800_n597# a_26_n597#
X0 a_325_n500# a_262_n597# a_207_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X1 a_561_n500# a_498_n597# a_443_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X2 a_n265_n500# a_n328_n597# a_n383_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X3 a_797_n500# a_734_n597# a_679_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X4 a_89_n500# a_26_n597# a_n29_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X5 a_207_n500# a_144_n597# a_89_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X6 a_n501_n500# a_n564_n597# a_n619_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X7 a_n147_n500# a_n210_n597# a_n265_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=300000u
X8 a_679_n500# a_616_n597# a_561_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X9 a_n737_n500# a_n800_n597# a_n855_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X10 a_443_n500# a_380_n597# a_325_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X11 a_n383_n500# a_n446_n597# a_n501_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X12 a_n619_n500# a_n682_n597# a_n737_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X13 a_n29_n500# a_n92_n597# a_n147_n500# w_n993_n719# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
.ends

.subckt sky130_fd_pr__nfet_01v8_Z85A38 a_1261_n500# a_n1319_n500# a_1577_n526# a_n287_n500#
+ a_n1061_n500# a_745_n500# a_29_n526# a_n1777_n526# a_n745_n526# a_1777_n500# a_n2351_n500#
+ a_803_n526# a_n2035_n526# a_229_n500# a_n1577_n500# a_2035_n500# a_1835_n526# a_n229_n526#
+ a_n545_n500# a_287_n526# a_n1003_n526# a_2093_n526# a_1003_n500# a_1319_n526# a_n2293_n526#
+ a_1061_n526# a_n29_n500# a_487_n500# a_2293_n500# a_n1835_n500# a_n1519_n526# a_n487_n526#
+ a_n1261_n526# a_1519_n500# a_n803_n500# a_545_n526# a_n2093_n500# VSUBS
X0 a_n1577_n500# a_n1777_n526# a_n1835_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X1 a_1519_n500# a_1319_n526# a_1261_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X2 a_n1061_n500# a_n1261_n526# a_n1319_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X3 a_1003_n500# a_803_n526# a_745_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X4 a_487_n500# a_287_n526# a_229_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X5 a_745_n500# a_545_n526# a_487_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X6 a_2035_n500# a_1835_n526# a_1777_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X7 a_1777_n500# a_1577_n526# a_1519_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 a_1261_n500# a_1061_n526# a_1003_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X9 a_n1835_n500# a_n2035_n526# a_n2093_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X10 a_n2093_n500# a_n2293_n526# a_n2351_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X11 a_n29_n500# a_n229_n526# a_n287_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X12 a_229_n500# a_29_n526# a_n29_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X13 a_n1319_n500# a_n1519_n526# a_n1577_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X14 a_n545_n500# a_n745_n526# a_n803_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X15 a_2293_n500# a_2093_n526# a_2035_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X16 a_n803_n500# a_n1003_n526# a_n1061_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X17 a_n287_n500# a_n487_n526# a_n545_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_U3DWQW a_n345_n800# a_129_n800# a_n503_n800# a_29_n826#
+ a_n661_n800# a_n129_n826# a_287_n800# a_187_n826# a_n287_n826# a_445_n800# a_345_n826#
+ a_n445_n826# a_603_n800# a_503_n826# a_n603_n826# a_761_n800# a_661_n826# a_n29_n800#
+ a_n761_n826# a_n187_n800# a_n819_n800# VSUBS
X0 a_n661_n800# a_n761_n826# a_n819_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X1 a_n187_n800# a_n287_n826# a_n345_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X2 a_761_n800# a_661_n826# a_603_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X3 a_287_n800# a_187_n826# a_129_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X4 a_n345_n800# a_n445_n826# a_n503_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X5 a_129_n800# a_29_n826# a_n29_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X6 a_445_n800# a_345_n826# a_287_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=500000u
X7 a_n503_n800# a_n603_n826# a_n661_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X8 a_n29_n800# a_n129_n826# a_n187_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X9 a_603_n800# a_503_n826# a_445_n800# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_2J7QF2 a_147_n526# a_n501_n500# a_561_n500# a_n383_n500#
+ a_29_n526# a_n737_n500# a_n561_n526# a_443_n500# a_n265_n500# a_n443_n526# a_n619_n500#
+ a_325_n500# a_501_n526# a_679_n500# a_n147_n500# a_n325_n526# a_383_n526# a_n679_n526#
+ a_207_n500# a_n29_n500# a_n207_n526# a_265_n526# a_619_n526# a_89_n500# a_n89_n526#
+ VSUBS
X0 a_n383_n500# a_n443_n526# a_n501_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X1 a_n619_n500# a_n679_n526# a_n737_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X2 a_n29_n500# a_n89_n526# a_n147_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X3 a_325_n500# a_265_n526# a_207_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X4 a_n265_n500# a_n325_n526# a_n383_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=300000u
X5 a_561_n500# a_501_n526# a_443_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=300000u
X6 a_89_n500# a_29_n526# a_n29_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=300000u
X7 a_207_n500# a_147_n526# a_89_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X8 a_n501_n500# a_n561_n526# a_n619_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X9 a_n147_n500# a_n207_n526# a_n265_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
X10 a_679_n500# a_619_n526# a_561_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=300000u
X11 a_443_n500# a_383_n526# a_325_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=300000u
.ends

.subckt opamp POS NEG VSS VDD EA_OUT BIAS_CUR
Xsky130_fd_pr__nfet_01v8_lvt_A3UXRA_0 VSS VSS VSS P1 VSS VSS VSS P1 VSS VSS P1 VSS
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS P1 VSS
+ VSS VSS P1 VSS P1 VSS VSS VSS P1 VSS VSS P1 VSS P1 P1 P1 VSS P1 VSS P1 VSS VSS P1
+ VSS VSS VSS P1 P1 P1 VSS VSS VSS VSS P1 VSS VSS P1 P1 VSS VSS VSS VSS VSS P1 VSS
+ P1 VSS VSS P1 VSS P1 P1 P1 VSS VSS P1 P1 VSS VSS VSS VSS VSS P1 P1 VSS VSS VSS VSS
+ VSS VSS VSS P1 P1 VSS VSS VSS VSS VSS VSS VSS P1 VSS P1 VSS VSS VSS VSS VSS VSS
+ P1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS P1 VSS P1 VSS
+ VSS VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS P1 VSS
+ VSS VSS VSS VSS VSS P1 VSS P1 VSS VSS VSS P1 VSS VSS VSS VSS VSS P1 VSS VSS VSS
+ P1 VSS P1 VSS VSS P1 P1 VSS VSS VSS P1 VSS VSS VSS VSS P1 P1 P1 VSS P1 P1 VSS VSS
+ P1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS P1 VSS VSS P1
+ VSS P1 P1 VSS P1 VSS P1 P1 P1 VSS VSS VSS P1 VSS VSS VSS VSS P1 VSS P1 VSS VSS P1
+ VSS VSS P1 VSS P1 VSS VSS P1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS
+ VSS VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS VSS VSS VSS P1 VSS P1 VSS VSS P1 VSS VSS
+ VSS VSS VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS P1 VSS P1 VSS P1 VSS VSS VSS VSS VSS
+ VSS P1 VSS VSS VSS VSS VSS P1 VSS P1 VSS P1 VSS VSS VSS VSS VSS VSS P1 VSS P1 VSS
+ VSS VSS P1 VSS VSS P1 VSS P1 VSS VSS VSS P1 VSS VSS VSS VSS VSS P1 VSS P1 VSS P1
+ VSS VSS VSS P1 VSS P1 VSS VSS P1 VSS VSS VSS P1 P1 VSS P1 P1 VSS VSS P1 VSS VSS
+ VSS VSS P1 P1 VSS VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS VSS P1 P1 VSS VSS VSS P1
+ VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS VSS VSS
+ VSS P1 VSS P1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS
+ P1 VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS
+ VSS VSS VSS VSS P1 VSS VSS P1 VSS VSS P1 VSS VSS VSS VSS VSS VSS VSS P1 P1 VSS VSS
+ VSS VSS VSS VSS P1 VSS VSS VSS P1 VSS P1 P1 P1 P1 VSS VSS VSS VSS P1 VSS P1 VSS
+ VSS VSS VSS VSS VSS VSS P1 VSS P1 VSS VSS VSS VSS VSS P1 VSS P1 VSS VSS VSS VSS
+ P1 P1 P1 VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS P1 VSS VSS VSS VSS
+ P1 VSS VSS P1 VSS VSS VSS VSS VSS VSS P1 P1 VSS VSS VSS P1 VSS VSS VSS VSS VSS VSS
+ P1 VSS VSS VSS VSS P1 VSS sky130_fd_pr__nfet_01v8_lvt_A3UXRA
Xsky130_fd_pr__pfet_01v8_477Z4B_0 NEG_D NEG_2 VDD VDD VDD NEG_D NEG_D NEG_D VDD NEG_2
+ NEG_D NEG_D NEG_D NEG_D VDD VDD VDD NEG_D VDD NEG_D NEG_D NEG_D VDD NEG_D NEG_D
+ NEG_D NEG_2 VDD VDD NEG_D sky130_fd_pr__pfet_01v8_477Z4B
Xsky130_fd_pr__pfet_01v8_477Z4B_1 POS_D EA_OUT VDD VDD VDD POS_D POS_D POS_D VDD EA_OUT
+ POS_D POS_D POS_D POS_D VDD VDD VDD POS_D VDD POS_D POS_D POS_D VDD POS_D POS_D
+ POS_D EA_OUT VDD VDD POS_D sky130_fd_pr__pfet_01v8_477Z4B
Xsky130_fd_pr__nfet_01v8_Z85A38_0 VSS VSS BIAS_CUR VSS P1 VSS BIAS_CUR BIAS_CUR BIAS_CUR
+ VSS VSS BIAS_CUR BIAS_CUR VSS BIAS_CUR P1 BIAS_CUR BIAS_CUR BIAS_CUR BIAS_CUR BIAS_CUR
+ VSS P1 BIAS_CUR VSS BIAS_CUR P1 BIAS_CUR VSS VSS BIAS_CUR BIAS_CUR BIAS_CUR BIAS_CUR
+ VSS BIAS_CUR P1 VSS sky130_fd_pr__nfet_01v8_Z85A38
Xsky130_fd_pr__nfet_01v8_U3DWQW_0 POS_D P1 P1 NEG NEG_D NEG POS_D POS POS P1 POS POS
+ NEG_D NEG NEG P1 P1 NEG_D P1 P1 P1 VSS sky130_fd_pr__nfet_01v8_U3DWQW
Xsky130_fd_pr__nfet_01v8_2J7QF2_0 NEG_2 VSS EA_OUT EA_OUT NEG_2 VSS NEG_2 VSS VSS
+ NEG_2 NEG_2 NEG_2 NEG_2 VSS NEG_2 NEG_2 NEG_2 NEG_2 VSS VSS NEG_2 NEG_2 NEG_2 EA_OUT
+ NEG_2 VSS sky130_fd_pr__nfet_01v8_2J7QF2
.ends

.subckt ulqc_ldo VIN VSS ADJ BGR_IN EA_OUT OUT
Xpower_transistor_0 VIN EA_OUT opamp_0/BIAS_CUR OUT power_transistor
Xopamp_0 ADJ BGR_IN VSS VIN EA_OUT opamp_0/BIAS_CUR opamp
.ends

.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2
+ wb_clk_i wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i[3] wbs_sel_i[2] wbs_sel_i[1]
+ wbs_sel_i[0] wbs_dat_i[31] wbs_dat_i[30] wbs_dat_i[29] wbs_dat_i[28] wbs_dat_i[27]
+ wbs_dat_i[26] wbs_dat_i[25] wbs_dat_i[24] wbs_dat_i[23] wbs_dat_i[22] wbs_dat_i[21]
+ wbs_dat_i[20] wbs_dat_i[19] wbs_dat_i[18] wbs_dat_i[17] wbs_dat_i[16] wbs_dat_i[15]
+ wbs_dat_i[14] wbs_dat_i[13] wbs_dat_i[12] wbs_dat_i[11] wbs_dat_i[10] wbs_dat_i[9]
+ wbs_dat_i[8] wbs_dat_i[7] wbs_dat_i[6] wbs_dat_i[5] wbs_dat_i[4] wbs_dat_i[3] wbs_dat_i[2]
+ wbs_dat_i[1] wbs_dat_i[0] wbs_adr_i[31] wbs_adr_i[30] wbs_adr_i[29] wbs_adr_i[28]
+ wbs_adr_i[27] wbs_adr_i[26] wbs_adr_i[25] wbs_adr_i[24] wbs_adr_i[23] wbs_adr_i[22]
+ wbs_adr_i[21] wbs_adr_i[20] wbs_adr_i[19] wbs_adr_i[18] wbs_adr_i[17] wbs_adr_i[16]
+ wbs_adr_i[15] wbs_adr_i[14] wbs_adr_i[13] wbs_adr_i[12] wbs_adr_i[11] wbs_adr_i[10]
+ wbs_adr_i[9] wbs_adr_i[8] wbs_adr_i[7] wbs_adr_i[6] wbs_adr_i[5] wbs_adr_i[4] wbs_adr_i[3]
+ wbs_adr_i[2] wbs_adr_i[1] wbs_adr_i[0] wbs_ack_o wbs_dat_o[31] wbs_dat_o[30] wbs_dat_o[29]
+ wbs_dat_o[28] wbs_dat_o[27] wbs_dat_o[26] wbs_dat_o[25] wbs_dat_o[24] wbs_dat_o[23]
+ wbs_dat_o[22] wbs_dat_o[21] wbs_dat_o[20] wbs_dat_o[19] wbs_dat_o[18] wbs_dat_o[17]
+ wbs_dat_o[16] wbs_dat_o[15] wbs_dat_o[14] wbs_dat_o[13] wbs_dat_o[12] wbs_dat_o[11]
+ wbs_dat_o[10] wbs_dat_o[9] wbs_dat_o[8] wbs_dat_o[7] wbs_dat_o[6] wbs_dat_o[5] wbs_dat_o[4]
+ wbs_dat_o[3] wbs_dat_o[2] wbs_dat_o[1] wbs_dat_o[0] la_data_in[127] la_data_in[126]
+ la_data_in[125] la_data_in[124] la_data_in[123] la_data_in[122] la_data_in[121]
+ la_data_in[120] la_data_in[119] la_data_in[118] la_data_in[117] la_data_in[116]
+ la_data_in[115] la_data_in[114] la_data_in[113] la_data_in[112] la_data_in[111]
+ la_data_in[110] la_data_in[109] la_data_in[108] la_data_in[107] la_data_in[106]
+ la_data_in[105] la_data_in[104] la_data_in[103] la_data_in[102] la_data_in[101]
+ la_data_in[100] la_data_in[99] la_data_in[98] la_data_in[97] la_data_in[96] la_data_in[95]
+ la_data_in[94] la_data_in[93] la_data_in[92] la_data_in[91] la_data_in[90] la_data_in[89]
+ la_data_in[88] la_data_in[87] la_data_in[86] la_data_in[85] la_data_in[84] la_data_in[83]
+ la_data_in[82] la_data_in[81] la_data_in[80] la_data_in[79] la_data_in[78] la_data_in[77]
+ la_data_in[76] la_data_in[75] la_data_in[74] la_data_in[73] la_data_in[72] la_data_in[71]
+ la_data_in[70] la_data_in[69] la_data_in[68] la_data_in[67] la_data_in[66] la_data_in[65]
+ la_data_in[64] la_data_in[63] la_data_in[62] la_data_in[61] la_data_in[60] la_data_in[59]
+ la_data_in[58] la_data_in[57] la_data_in[56] la_data_in[55] la_data_in[54] la_data_in[53]
+ la_data_in[52] la_data_in[51] la_data_in[50] la_data_in[49] la_data_in[48] la_data_in[47]
+ la_data_in[46] la_data_in[45] la_data_in[44] la_data_in[43] la_data_in[42] la_data_in[41]
+ la_data_in[40] la_data_in[39] la_data_in[38] la_data_in[37] la_data_in[36] la_data_in[35]
+ la_data_in[34] la_data_in[33] la_data_in[32] la_data_in[31] la_data_in[30] la_data_in[29]
+ la_data_in[28] la_data_in[27] la_data_in[26] la_data_in[25] la_data_in[24] la_data_in[23]
+ la_data_in[22] la_data_in[21] la_data_in[20] la_data_in[19] la_data_in[18] la_data_in[17]
+ la_data_in[16] la_data_in[15] la_data_in[14] la_data_in[13] la_data_in[12] la_data_in[11]
+ la_data_in[10] la_data_in[9] la_data_in[8] la_data_in[7] la_data_in[6] la_data_in[5]
+ la_data_in[4] la_data_in[3] la_data_in[2] la_data_in[1] la_data_in[0] la_data_out[127]
+ la_data_out[126] la_data_out[125] la_data_out[124] la_data_out[123] la_data_out[122]
+ la_data_out[121] la_data_out[120] la_data_out[119] la_data_out[118] la_data_out[117]
+ la_data_out[116] la_data_out[115] la_data_out[114] la_data_out[113] la_data_out[112]
+ la_data_out[111] la_data_out[110] la_data_out[109] la_data_out[108] la_data_out[107]
+ la_data_out[106] la_data_out[105] la_data_out[104] la_data_out[103] la_data_out[102]
+ la_data_out[101] la_data_out[100] la_data_out[99] la_data_out[98] la_data_out[97]
+ la_data_out[96] la_data_out[95] la_data_out[94] la_data_out[93] la_data_out[92]
+ la_data_out[91] la_data_out[90] la_data_out[89] la_data_out[88] la_data_out[87]
+ la_data_out[86] la_data_out[85] la_data_out[84] la_data_out[83] la_data_out[82]
+ la_data_out[81] la_data_out[80] la_data_out[79] la_data_out[78] la_data_out[77]
+ la_data_out[76] la_data_out[75] la_data_out[74] la_data_out[73] la_data_out[72]
+ la_data_out[71] la_data_out[70] la_data_out[69] la_data_out[68] la_data_out[67]
+ la_data_out[66] la_data_out[65] la_data_out[64] la_data_out[63] la_data_out[62]
+ la_data_out[61] la_data_out[60] la_data_out[59] la_data_out[58] la_data_out[57]
+ la_data_out[56] la_data_out[55] la_data_out[54] la_data_out[53] la_data_out[52]
+ la_data_out[51] la_data_out[50] la_data_out[49] la_data_out[48] la_data_out[47]
+ la_data_out[46] la_data_out[45] la_data_out[44] la_data_out[43] la_data_out[42]
+ la_data_out[41] la_data_out[40] la_data_out[39] la_data_out[38] la_data_out[37]
+ la_data_out[36] la_data_out[35] la_data_out[34] la_data_out[33] la_data_out[32]
+ la_data_out[31] la_data_out[30] la_data_out[29] la_data_out[28] la_data_out[27]
+ la_data_out[26] la_data_out[25] la_data_out[24] la_data_out[23] la_data_out[22]
+ la_data_out[21] la_data_out[20] la_data_out[19] la_data_out[18] la_data_out[17]
+ la_data_out[16] la_data_out[15] la_data_out[14] la_data_out[13] la_data_out[12]
+ la_data_out[11] la_data_out[10] la_data_out[9] la_data_out[8] la_data_out[7] la_data_out[6]
+ la_data_out[5] la_data_out[4] la_data_out[3] la_data_out[2] la_data_out[1] la_data_out[0]
+ io_in[26] io_in[25] io_in[24] io_in[23] io_in[22] io_in[21] io_in[20] io_in[19]
+ io_in[18] io_in[17] io_in[16] io_in[15] io_in[14] io_in[13] io_in[12] io_in[11]
+ io_in[10] io_in[9] io_in[8] io_in[7] io_in[6] io_in[5] io_in[4] io_in[3] io_in[2]
+ io_in[1] io_in[0] io_in_3v3[26] io_in_3v3[25] io_in_3v3[24] io_in_3v3[23] io_in_3v3[22]
+ io_in_3v3[21] io_in_3v3[20] io_in_3v3[19] io_in_3v3[18] io_in_3v3[17] io_in_3v3[16]
+ io_in_3v3[15] io_in_3v3[14] io_in_3v3[13] io_in_3v3[12] io_in_3v3[11] io_in_3v3[10]
+ io_in_3v3[9] io_in_3v3[8] io_in_3v3[7] io_in_3v3[6] io_in_3v3[5] io_in_3v3[4] io_in_3v3[3]
+ io_in_3v3[2] io_in_3v3[1] io_in_3v3[0] user_clock2 io_out[26] io_out[25] io_out[24]
+ io_out[23] io_out[22] io_out[21] io_out[20] io_out[19] io_out[18] io_out[17] io_out[16]
+ io_out[15] io_out[14] io_out[13] io_out[12] io_out[11] io_out[10] io_out[9] io_out[8]
+ io_out[7] io_out[6] io_out[5] io_out[4] io_out[3] io_out[2] io_out[1] io_out[0]
+ io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22] io_oeb[21] io_oeb[20] io_oeb[19]
+ io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15] io_oeb[14] io_oeb[13] io_oeb[12] io_oeb[11]
+ io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[7] io_oeb[6] io_oeb[5] io_oeb[4] io_oeb[3]
+ io_oeb[2] io_oeb[1] io_oeb[0] gpio_analog[17] gpio_analog[16] gpio_analog[15] gpio_analog[14]
+ gpio_analog[13] gpio_analog[12] gpio_analog[11] gpio_analog[10] gpio_analog[9] gpio_analog[8]
+ gpio_analog[7] gpio_analog[6] gpio_analog[5] gpio_analog[4] gpio_analog[3] gpio_analog[2]
+ gpio_analog[1] gpio_analog[0] gpio_noesd[17] gpio_noesd[16] gpio_noesd[15] gpio_noesd[14]
+ gpio_noesd[13] gpio_noesd[12] gpio_noesd[11] gpio_noesd[10] gpio_noesd[9] gpio_noesd[8]
+ gpio_noesd[7] gpio_noesd[6] gpio_noesd[5] gpio_noesd[4] gpio_noesd[3] gpio_noesd[2]
+ gpio_noesd[1] gpio_noesd[0] io_analog[10] io_analog[9] io_analog[8] io_analog[7]
+ io_analog[6] io_analog[5] io_analog[4] io_analog[3] io_analog[2] io_analog[1] io_analog[0]
+ io_clamp_high[2] io_clamp_high[1] io_clamp_high[0] io_clamp_low[2] io_clamp_low[1]
+ io_clamp_low[0] user_irq[2] user_irq[1] user_irq[0] la_oenb[127] la_oenb[126] la_oenb[125]
+ la_oenb[124] la_oenb[123] la_oenb[122] la_oenb[121] la_oenb[120] la_oenb[119] la_oenb[118]
+ la_oenb[117] la_oenb[116] la_oenb[115] la_oenb[114] la_oenb[113] la_oenb[112] la_oenb[111]
+ la_oenb[110] la_oenb[109] la_oenb[108] la_oenb[107] la_oenb[106] la_oenb[105] la_oenb[104]
+ la_oenb[103] la_oenb[102] la_oenb[101] la_oenb[100] la_oenb[99] la_oenb[98] la_oenb[97]
+ la_oenb[96] la_oenb[95] la_oenb[94] la_oenb[93] la_oenb[92] la_oenb[91] la_oenb[90]
+ la_oenb[89] la_oenb[88] la_oenb[87] la_oenb[86] la_oenb[85] la_oenb[84] la_oenb[83]
+ la_oenb[82] la_oenb[81] la_oenb[80] la_oenb[79] la_oenb[78] la_oenb[77] la_oenb[76]
+ la_oenb[75] la_oenb[74] la_oenb[73] la_oenb[72] la_oenb[71] la_oenb[70] la_oenb[69]
+ la_oenb[68] la_oenb[67] la_oenb[66] la_oenb[65] la_oenb[64] la_oenb[63] la_oenb[62]
+ la_oenb[61] la_oenb[60] la_oenb[59] la_oenb[58] la_oenb[57] la_oenb[56] la_oenb[55]
+ la_oenb[54] la_oenb[53] la_oenb[52] la_oenb[51] la_oenb[50] la_oenb[49] la_oenb[48]
+ la_oenb[47] la_oenb[46] la_oenb[45] la_oenb[44] la_oenb[43] la_oenb[42] la_oenb[41]
+ la_oenb[40] la_oenb[39] la_oenb[38] la_oenb[37] la_oenb[36] la_oenb[35] la_oenb[34]
+ la_oenb[33] la_oenb[32] la_oenb[31] la_oenb[30] la_oenb[29] la_oenb[28] la_oenb[27]
+ la_oenb[26] la_oenb[25] la_oenb[24] la_oenb[23] la_oenb[22] la_oenb[21] la_oenb[20]
+ la_oenb[19] la_oenb[18] la_oenb[17] la_oenb[16] la_oenb[15] la_oenb[14] la_oenb[13]
+ la_oenb[12] la_oenb[11] la_oenb[10] la_oenb[9] la_oenb[8] la_oenb[7] la_oenb[6]
+ la_oenb[5] la_oenb[4] la_oenb[3] la_oenb[2] la_oenb[1] la_oenb[0]
Xulqc_ldo_0 io_analog[4] vssa1 io_analog[3] io_analog[7] io_analog[2] io_analog[0]
+ ulqc_ldo
.ends

