magic
tech sky130A
magscale 1 2
timestamp 1697794388
<< error_p >>
rect -623 572 -565 578
rect -407 572 -349 578
rect -191 572 -133 578
rect 25 572 83 578
rect 241 572 299 578
rect 457 572 515 578
rect 673 572 731 578
rect -623 538 -611 572
rect -407 538 -395 572
rect -191 538 -179 572
rect 25 538 37 572
rect 241 538 253 572
rect 457 538 469 572
rect 673 538 685 572
rect -623 532 -565 538
rect -407 532 -349 538
rect -191 532 -133 538
rect 25 532 83 538
rect 241 532 299 538
rect 457 532 515 538
rect 673 532 731 538
rect -731 -538 -673 -532
rect -515 -538 -457 -532
rect -299 -538 -241 -532
rect -83 -538 -25 -532
rect 133 -538 191 -532
rect 349 -538 407 -532
rect 565 -538 623 -532
rect -731 -572 -719 -538
rect -515 -572 -503 -538
rect -299 -572 -287 -538
rect -83 -572 -71 -538
rect 133 -572 145 -538
rect 349 -572 361 -538
rect 565 -572 577 -538
rect -731 -578 -673 -572
rect -515 -578 -457 -572
rect -299 -578 -241 -572
rect -83 -578 -25 -572
rect 133 -578 191 -572
rect 349 -578 407 -572
rect 565 -578 623 -572
<< nmos >>
rect -727 -500 -677 500
rect -619 -500 -569 500
rect -511 -500 -461 500
rect -403 -500 -353 500
rect -295 -500 -245 500
rect -187 -500 -137 500
rect -79 -500 -29 500
rect 29 -500 79 500
rect 137 -500 187 500
rect 245 -500 295 500
rect 353 -500 403 500
rect 461 -500 511 500
rect 569 -500 619 500
rect 677 -500 727 500
<< ndiff >>
rect -785 488 -727 500
rect -785 -488 -773 488
rect -739 -488 -727 488
rect -785 -500 -727 -488
rect -677 488 -619 500
rect -677 -488 -665 488
rect -631 -488 -619 488
rect -677 -500 -619 -488
rect -569 488 -511 500
rect -569 -488 -557 488
rect -523 -488 -511 488
rect -569 -500 -511 -488
rect -461 488 -403 500
rect -461 -488 -449 488
rect -415 -488 -403 488
rect -461 -500 -403 -488
rect -353 488 -295 500
rect -353 -488 -341 488
rect -307 -488 -295 488
rect -353 -500 -295 -488
rect -245 488 -187 500
rect -245 -488 -233 488
rect -199 -488 -187 488
rect -245 -500 -187 -488
rect -137 488 -79 500
rect -137 -488 -125 488
rect -91 -488 -79 488
rect -137 -500 -79 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 79 488 137 500
rect 79 -488 91 488
rect 125 -488 137 488
rect 79 -500 137 -488
rect 187 488 245 500
rect 187 -488 199 488
rect 233 -488 245 488
rect 187 -500 245 -488
rect 295 488 353 500
rect 295 -488 307 488
rect 341 -488 353 488
rect 295 -500 353 -488
rect 403 488 461 500
rect 403 -488 415 488
rect 449 -488 461 488
rect 403 -500 461 -488
rect 511 488 569 500
rect 511 -488 523 488
rect 557 -488 569 488
rect 511 -500 569 -488
rect 619 488 677 500
rect 619 -488 631 488
rect 665 -488 677 488
rect 619 -500 677 -488
rect 727 488 785 500
rect 727 -488 739 488
rect 773 -488 785 488
rect 727 -500 785 -488
<< ndiffc >>
rect -773 -488 -739 488
rect -665 -488 -631 488
rect -557 -488 -523 488
rect -449 -488 -415 488
rect -341 -488 -307 488
rect -233 -488 -199 488
rect -125 -488 -91 488
rect -17 -488 17 488
rect 91 -488 125 488
rect 199 -488 233 488
rect 307 -488 341 488
rect 415 -488 449 488
rect 523 -488 557 488
rect 631 -488 665 488
rect 739 -488 773 488
<< poly >>
rect -627 572 -561 588
rect -627 538 -611 572
rect -577 538 -561 572
rect -727 500 -677 526
rect -627 522 -561 538
rect -411 572 -345 588
rect -411 538 -395 572
rect -361 538 -345 572
rect -619 500 -569 522
rect -511 500 -461 526
rect -411 522 -345 538
rect -195 572 -129 588
rect -195 538 -179 572
rect -145 538 -129 572
rect -403 500 -353 522
rect -295 500 -245 526
rect -195 522 -129 538
rect 21 572 87 588
rect 21 538 37 572
rect 71 538 87 572
rect -187 500 -137 522
rect -79 500 -29 526
rect 21 522 87 538
rect 237 572 303 588
rect 237 538 253 572
rect 287 538 303 572
rect 29 500 79 522
rect 137 500 187 526
rect 237 522 303 538
rect 453 572 519 588
rect 453 538 469 572
rect 503 538 519 572
rect 245 500 295 522
rect 353 500 403 526
rect 453 522 519 538
rect 669 572 735 588
rect 669 538 685 572
rect 719 538 735 572
rect 461 500 511 522
rect 569 500 619 526
rect 669 522 735 538
rect 677 500 727 522
rect -727 -522 -677 -500
rect -735 -538 -669 -522
rect -619 -526 -569 -500
rect -511 -522 -461 -500
rect -735 -572 -719 -538
rect -685 -572 -669 -538
rect -735 -588 -669 -572
rect -519 -538 -453 -522
rect -403 -526 -353 -500
rect -295 -522 -245 -500
rect -519 -572 -503 -538
rect -469 -572 -453 -538
rect -519 -588 -453 -572
rect -303 -538 -237 -522
rect -187 -526 -137 -500
rect -79 -522 -29 -500
rect -303 -572 -287 -538
rect -253 -572 -237 -538
rect -303 -588 -237 -572
rect -87 -538 -21 -522
rect 29 -526 79 -500
rect 137 -522 187 -500
rect -87 -572 -71 -538
rect -37 -572 -21 -538
rect -87 -588 -21 -572
rect 129 -538 195 -522
rect 245 -526 295 -500
rect 353 -522 403 -500
rect 129 -572 145 -538
rect 179 -572 195 -538
rect 129 -588 195 -572
rect 345 -538 411 -522
rect 461 -526 511 -500
rect 569 -522 619 -500
rect 345 -572 361 -538
rect 395 -572 411 -538
rect 345 -588 411 -572
rect 561 -538 627 -522
rect 677 -526 727 -500
rect 561 -572 577 -538
rect 611 -572 627 -538
rect 561 -588 627 -572
<< polycont >>
rect -611 538 -577 572
rect -395 538 -361 572
rect -179 538 -145 572
rect 37 538 71 572
rect 253 538 287 572
rect 469 538 503 572
rect 685 538 719 572
rect -719 -572 -685 -538
rect -503 -572 -469 -538
rect -287 -572 -253 -538
rect -71 -572 -37 -538
rect 145 -572 179 -538
rect 361 -572 395 -538
rect 577 -572 611 -538
<< locali >>
rect -627 538 -611 572
rect -577 538 -561 572
rect -411 538 -395 572
rect -361 538 -345 572
rect -195 538 -179 572
rect -145 538 -129 572
rect 21 538 37 572
rect 71 538 87 572
rect 237 538 253 572
rect 287 538 303 572
rect 453 538 469 572
rect 503 538 519 572
rect 669 538 685 572
rect 719 538 735 572
rect -773 488 -739 504
rect -773 -504 -739 -488
rect -665 488 -631 504
rect -665 -504 -631 -488
rect -557 488 -523 504
rect -557 -504 -523 -488
rect -449 488 -415 504
rect -449 -504 -415 -488
rect -341 488 -307 504
rect -341 -504 -307 -488
rect -233 488 -199 504
rect -233 -504 -199 -488
rect -125 488 -91 504
rect -125 -504 -91 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 91 488 125 504
rect 91 -504 125 -488
rect 199 488 233 504
rect 199 -504 233 -488
rect 307 488 341 504
rect 307 -504 341 -488
rect 415 488 449 504
rect 415 -504 449 -488
rect 523 488 557 504
rect 523 -504 557 -488
rect 631 488 665 504
rect 631 -504 665 -488
rect 739 488 773 504
rect 739 -504 773 -488
rect -735 -572 -719 -538
rect -685 -572 -669 -538
rect -519 -572 -503 -538
rect -469 -572 -453 -538
rect -303 -572 -287 -538
rect -253 -572 -237 -538
rect -87 -572 -71 -538
rect -37 -572 -21 -538
rect 129 -572 145 -538
rect 179 -572 195 -538
rect 345 -572 361 -538
rect 395 -572 411 -538
rect 561 -572 577 -538
rect 611 -572 627 -538
<< viali >>
rect -611 538 -577 572
rect -395 538 -361 572
rect -179 538 -145 572
rect 37 538 71 572
rect 253 538 287 572
rect 469 538 503 572
rect 685 538 719 572
rect -773 -488 -739 488
rect -665 -488 -631 488
rect -557 -488 -523 488
rect -449 -488 -415 488
rect -341 -488 -307 488
rect -233 -488 -199 488
rect -125 -488 -91 488
rect -17 -488 17 488
rect 91 -488 125 488
rect 199 -488 233 488
rect 307 -488 341 488
rect 415 -488 449 488
rect 523 -488 557 488
rect 631 -488 665 488
rect 739 -488 773 488
rect -719 -572 -685 -538
rect -503 -572 -469 -538
rect -287 -572 -253 -538
rect -71 -572 -37 -538
rect 145 -572 179 -538
rect 361 -572 395 -538
rect 577 -572 611 -538
<< metal1 >>
rect -623 572 -565 578
rect -623 538 -611 572
rect -577 538 -565 572
rect -623 532 -565 538
rect -407 572 -349 578
rect -407 538 -395 572
rect -361 538 -349 572
rect -407 532 -349 538
rect -191 572 -133 578
rect -191 538 -179 572
rect -145 538 -133 572
rect -191 532 -133 538
rect 25 572 83 578
rect 25 538 37 572
rect 71 538 83 572
rect 25 532 83 538
rect 241 572 299 578
rect 241 538 253 572
rect 287 538 299 572
rect 241 532 299 538
rect 457 572 515 578
rect 457 538 469 572
rect 503 538 515 572
rect 457 532 515 538
rect 673 572 731 578
rect 673 538 685 572
rect 719 538 731 572
rect 673 532 731 538
rect -779 488 -733 500
rect -779 -488 -773 488
rect -739 -488 -733 488
rect -779 -500 -733 -488
rect -671 488 -625 500
rect -671 -488 -665 488
rect -631 -488 -625 488
rect -671 -500 -625 -488
rect -563 488 -517 500
rect -563 -488 -557 488
rect -523 -488 -517 488
rect -563 -500 -517 -488
rect -455 488 -409 500
rect -455 -488 -449 488
rect -415 -488 -409 488
rect -455 -500 -409 -488
rect -347 488 -301 500
rect -347 -488 -341 488
rect -307 -488 -301 488
rect -347 -500 -301 -488
rect -239 488 -193 500
rect -239 -488 -233 488
rect -199 -488 -193 488
rect -239 -500 -193 -488
rect -131 488 -85 500
rect -131 -488 -125 488
rect -91 -488 -85 488
rect -131 -500 -85 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 85 488 131 500
rect 85 -488 91 488
rect 125 -488 131 488
rect 85 -500 131 -488
rect 193 488 239 500
rect 193 -488 199 488
rect 233 -488 239 488
rect 193 -500 239 -488
rect 301 488 347 500
rect 301 -488 307 488
rect 341 -488 347 488
rect 301 -500 347 -488
rect 409 488 455 500
rect 409 -488 415 488
rect 449 -488 455 488
rect 409 -500 455 -488
rect 517 488 563 500
rect 517 -488 523 488
rect 557 -488 563 488
rect 517 -500 563 -488
rect 625 488 671 500
rect 625 -488 631 488
rect 665 -488 671 488
rect 625 -500 671 -488
rect 733 488 779 500
rect 733 -488 739 488
rect 773 -488 779 488
rect 733 -500 779 -488
rect -731 -538 -673 -532
rect -731 -572 -719 -538
rect -685 -572 -673 -538
rect -731 -578 -673 -572
rect -515 -538 -457 -532
rect -515 -572 -503 -538
rect -469 -572 -457 -538
rect -515 -578 -457 -572
rect -299 -538 -241 -532
rect -299 -572 -287 -538
rect -253 -572 -241 -538
rect -299 -578 -241 -572
rect -83 -538 -25 -532
rect -83 -572 -71 -538
rect -37 -572 -25 -538
rect -83 -578 -25 -572
rect 133 -538 191 -532
rect 133 -572 145 -538
rect 179 -572 191 -538
rect 133 -578 191 -572
rect 349 -538 407 -532
rect 349 -572 361 -538
rect 395 -572 407 -538
rect 349 -578 407 -572
rect 565 -538 623 -532
rect 565 -572 577 -538
rect 611 -572 623 -538
rect 565 -578 623 -572
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.25 m 1 nf 14 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
