magic
tech sky130A
magscale 1 2
timestamp 1697794388
<< pwell >>
rect -483 -1010 483 1010
<< nmos >>
rect -287 -800 -187 800
rect -129 -800 -29 800
rect 29 -800 129 800
rect 187 -800 287 800
<< ndiff >>
rect -345 788 -287 800
rect -345 -788 -333 788
rect -299 -788 -287 788
rect -345 -800 -287 -788
rect -187 788 -129 800
rect -187 -788 -175 788
rect -141 -788 -129 788
rect -187 -800 -129 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 129 788 187 800
rect 129 -788 141 788
rect 175 -788 187 788
rect 129 -800 187 -788
rect 287 788 345 800
rect 287 -788 299 788
rect 333 -788 345 788
rect 287 -800 345 -788
<< ndiffc >>
rect -333 -788 -299 788
rect -175 -788 -141 788
rect -17 -788 17 788
rect 141 -788 175 788
rect 299 -788 333 788
<< psubdiff >>
rect -447 940 -351 974
rect 351 940 447 974
rect -447 878 -413 940
rect 413 878 447 940
rect -447 -940 -413 -878
rect 413 -940 447 -878
rect -447 -974 -351 -940
rect 351 -974 447 -940
<< psubdiffcont >>
rect -351 940 351 974
rect -447 -878 -413 878
rect 413 -878 447 878
rect -351 -974 351 -940
<< poly >>
rect -287 872 -187 888
rect -287 838 -271 872
rect -203 838 -187 872
rect -287 800 -187 838
rect -129 872 -29 888
rect -129 838 -113 872
rect -45 838 -29 872
rect -129 800 -29 838
rect 29 872 129 888
rect 29 838 45 872
rect 113 838 129 872
rect 29 800 129 838
rect 187 872 287 888
rect 187 838 203 872
rect 271 838 287 872
rect 187 800 287 838
rect -287 -838 -187 -800
rect -287 -872 -271 -838
rect -203 -872 -187 -838
rect -287 -888 -187 -872
rect -129 -838 -29 -800
rect -129 -872 -113 -838
rect -45 -872 -29 -838
rect -129 -888 -29 -872
rect 29 -838 129 -800
rect 29 -872 45 -838
rect 113 -872 129 -838
rect 29 -888 129 -872
rect 187 -838 287 -800
rect 187 -872 203 -838
rect 271 -872 287 -838
rect 187 -888 287 -872
<< polycont >>
rect -271 838 -203 872
rect -113 838 -45 872
rect 45 838 113 872
rect 203 838 271 872
rect -271 -872 -203 -838
rect -113 -872 -45 -838
rect 45 -872 113 -838
rect 203 -872 271 -838
<< locali >>
rect -447 940 -351 974
rect 351 940 447 974
rect -447 878 -413 940
rect 413 878 447 940
rect -287 838 -271 872
rect -203 838 -187 872
rect -129 838 -113 872
rect -45 838 -29 872
rect 29 838 45 872
rect 113 838 129 872
rect 187 838 203 872
rect 271 838 287 872
rect -333 788 -299 804
rect -333 -804 -299 -788
rect -175 788 -141 804
rect -175 -804 -141 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 141 788 175 804
rect 141 -804 175 -788
rect 299 788 333 804
rect 299 -804 333 -788
rect -287 -872 -271 -838
rect -203 -872 -187 -838
rect -129 -872 -113 -838
rect -45 -872 -29 -838
rect 29 -872 45 -838
rect 113 -872 129 -838
rect 187 -872 203 -838
rect 271 -872 287 -838
rect -447 -940 -413 -878
rect 413 -940 447 -878
rect -447 -974 -351 -940
rect 351 -974 447 -940
<< viali >>
rect -271 838 -203 872
rect -113 838 -45 872
rect 45 838 113 872
rect 203 838 271 872
rect -333 -788 -299 788
rect -175 -788 -141 788
rect -17 -788 17 788
rect 141 -788 175 788
rect 299 -788 333 788
rect -271 -872 -203 -838
rect -113 -872 -45 -838
rect 45 -872 113 -838
rect 203 -872 271 -838
<< metal1 >>
rect -283 872 -191 878
rect -283 838 -271 872
rect -203 838 -191 872
rect -283 832 -191 838
rect -125 872 -33 878
rect -125 838 -113 872
rect -45 838 -33 872
rect -125 832 -33 838
rect 33 872 125 878
rect 33 838 45 872
rect 113 838 125 872
rect 33 832 125 838
rect 191 872 283 878
rect 191 838 203 872
rect 271 838 283 872
rect 191 832 283 838
rect -339 788 -293 800
rect -339 -788 -333 788
rect -299 -788 -293 788
rect -339 -800 -293 -788
rect -181 788 -135 800
rect -181 -788 -175 788
rect -141 -788 -135 788
rect -181 -800 -135 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 135 788 181 800
rect 135 -788 141 788
rect 175 -788 181 788
rect 135 -800 181 -788
rect 293 788 339 800
rect 293 -788 299 788
rect 333 -788 339 788
rect 293 -800 339 -788
rect -283 -838 -191 -832
rect -283 -872 -271 -838
rect -203 -872 -191 -838
rect -283 -878 -191 -872
rect -125 -838 -33 -832
rect -125 -872 -113 -838
rect -45 -872 -33 -838
rect -125 -878 -33 -872
rect 33 -838 125 -832
rect 33 -872 45 -838
rect 113 -872 125 -838
rect 33 -878 125 -872
rect 191 -838 283 -832
rect 191 -872 203 -838
rect 271 -872 283 -838
rect 191 -878 283 -872
<< properties >>
string FIXED_BBOX -430 -957 430 957
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
