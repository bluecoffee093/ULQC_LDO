magic
tech sky130A
magscale 1 2
timestamp 1697926267
<< pwell >>
rect -201 -2498 201 2498
<< psubdiff >>
rect -165 2428 -69 2462
rect 69 2428 165 2462
rect -165 2366 -131 2428
rect 131 2366 165 2428
rect -165 -2428 -131 -2366
rect 131 -2428 165 -2366
rect -165 -2462 -69 -2428
rect 69 -2462 165 -2428
<< psubdiffcont >>
rect -69 2428 69 2462
rect -165 -2366 -131 2366
rect 131 -2366 165 2366
rect -69 -2462 69 -2428
<< xpolycontact >>
rect -35 1900 35 2332
rect -35 -2332 35 -1900
<< ppolyres >>
rect -35 -1900 35 1900
<< locali >>
rect -165 2428 -69 2462
rect 69 2428 165 2462
rect -165 2366 -131 2428
rect 131 2366 165 2428
rect -165 -2428 -131 -2366
rect 131 -2428 165 -2366
rect -165 -2462 -69 -2428
rect 69 -2462 165 -2428
<< viali >>
rect -19 1917 19 2314
rect -19 -2314 19 -1917
<< metal1 >>
rect -25 2314 25 2326
rect -25 1917 -19 2314
rect 19 1917 25 2314
rect -25 1905 25 1917
rect -25 -1917 25 -1905
rect -25 -2314 -19 -1917
rect 19 -2314 25 -1917
rect -25 -2326 25 -2314
<< res0p35 >>
rect -37 -1902 37 1902
<< properties >>
string FIXED_BBOX -148 -2445 148 2445
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 19.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 18.473k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
