magic
tech sky130A
magscale 1 2
timestamp 1697926267
<< pwell >>
rect -201 -1478 201 1478
<< psubdiff >>
rect -165 1408 -69 1442
rect 69 1408 165 1442
rect -165 1346 -131 1408
rect 131 1346 165 1408
rect -165 -1408 -131 -1346
rect 131 -1408 165 -1346
rect -165 -1442 -69 -1408
rect 69 -1442 165 -1408
<< psubdiffcont >>
rect -69 1408 69 1442
rect -165 -1346 -131 1346
rect 131 -1346 165 1346
rect -69 -1442 69 -1408
<< xpolycontact >>
rect -35 880 35 1312
rect -35 -1312 35 -880
<< ppolyres >>
rect -35 -880 35 880
<< locali >>
rect -165 1408 -69 1442
rect 69 1408 165 1442
rect -165 1346 -131 1408
rect 131 1346 165 1408
rect -165 -1408 -131 -1346
rect 131 -1408 165 -1346
rect -165 -1442 -69 -1408
rect 69 -1442 165 -1408
<< viali >>
rect -19 897 19 1294
rect -19 -1294 19 -897
<< metal1 >>
rect -25 1294 25 1306
rect -25 897 -19 1294
rect 19 897 25 1294
rect -25 885 25 897
rect -25 -897 25 -885
rect -25 -1294 -19 -897
rect 19 -1294 25 -897
rect -25 -1306 25 -1294
<< res0p35 >>
rect -37 -882 37 882
<< properties >>
string FIXED_BBOX -148 -1425 148 1425
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 8.8 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 9.153k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
