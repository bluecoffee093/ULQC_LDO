magic
tech sky130A
magscale 1 2
timestamp 1697794388
<< nmos >>
rect -679 -500 -619 500
rect -561 -500 -501 500
rect -443 -500 -383 500
rect -325 -500 -265 500
rect -207 -500 -147 500
rect -89 -500 -29 500
rect 29 -500 89 500
rect 147 -500 207 500
rect 265 -500 325 500
rect 383 -500 443 500
rect 501 -500 561 500
rect 619 -500 679 500
<< ndiff >>
rect -737 488 -679 500
rect -737 -488 -725 488
rect -691 -488 -679 488
rect -737 -500 -679 -488
rect -619 488 -561 500
rect -619 -488 -607 488
rect -573 -488 -561 488
rect -619 -500 -561 -488
rect -501 488 -443 500
rect -501 -488 -489 488
rect -455 -488 -443 488
rect -501 -500 -443 -488
rect -383 488 -325 500
rect -383 -488 -371 488
rect -337 -488 -325 488
rect -383 -500 -325 -488
rect -265 488 -207 500
rect -265 -488 -253 488
rect -219 -488 -207 488
rect -265 -500 -207 -488
rect -147 488 -89 500
rect -147 -488 -135 488
rect -101 -488 -89 488
rect -147 -500 -89 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 89 488 147 500
rect 89 -488 101 488
rect 135 -488 147 488
rect 89 -500 147 -488
rect 207 488 265 500
rect 207 -488 219 488
rect 253 -488 265 488
rect 207 -500 265 -488
rect 325 488 383 500
rect 325 -488 337 488
rect 371 -488 383 488
rect 325 -500 383 -488
rect 443 488 501 500
rect 443 -488 455 488
rect 489 -488 501 488
rect 443 -500 501 -488
rect 561 488 619 500
rect 561 -488 573 488
rect 607 -488 619 488
rect 561 -500 619 -488
rect 679 488 737 500
rect 679 -488 691 488
rect 725 -488 737 488
rect 679 -500 737 -488
<< ndiffc >>
rect -725 -488 -691 488
rect -607 -488 -573 488
rect -489 -488 -455 488
rect -371 -488 -337 488
rect -253 -488 -219 488
rect -135 -488 -101 488
rect -17 -488 17 488
rect 101 -488 135 488
rect 219 -488 253 488
rect 337 -488 371 488
rect 455 -488 489 488
rect 573 -488 607 488
rect 691 -488 725 488
<< poly >>
rect -679 500 -619 526
rect -561 500 -501 526
rect -443 500 -383 526
rect -325 500 -265 526
rect -207 500 -147 526
rect -89 500 -29 526
rect 29 500 89 526
rect 147 500 207 526
rect 265 500 325 526
rect 383 500 443 526
rect 501 500 561 526
rect 619 500 679 526
rect -679 -526 -619 -500
rect -561 -526 -501 -500
rect -443 -526 -383 -500
rect -325 -526 -265 -500
rect -207 -526 -147 -500
rect -89 -526 -29 -500
rect 29 -526 89 -500
rect 147 -526 207 -500
rect 265 -526 325 -500
rect 383 -526 443 -500
rect 501 -526 561 -500
rect 619 -526 679 -500
<< locali >>
rect -725 488 -691 504
rect -725 -504 -691 -488
rect -607 488 -573 504
rect -607 -504 -573 -488
rect -489 488 -455 504
rect -489 -504 -455 -488
rect -371 488 -337 504
rect -371 -504 -337 -488
rect -253 488 -219 504
rect -253 -504 -219 -488
rect -135 488 -101 504
rect -135 -504 -101 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 101 488 135 504
rect 101 -504 135 -488
rect 219 488 253 504
rect 219 -504 253 -488
rect 337 488 371 504
rect 337 -504 371 -488
rect 455 488 489 504
rect 455 -504 489 -488
rect 573 488 607 504
rect 573 -504 607 -488
rect 691 488 725 504
rect 691 -504 725 -488
<< viali >>
rect -725 -488 -691 488
rect -607 -488 -573 488
rect -489 -488 -455 488
rect -371 -488 -337 488
rect -253 -488 -219 488
rect -135 -488 -101 488
rect -17 -488 17 488
rect 101 -488 135 488
rect 219 -488 253 488
rect 337 -488 371 488
rect 455 -488 489 488
rect 573 -488 607 488
rect 691 -488 725 488
<< metal1 >>
rect -731 488 -685 500
rect -731 -488 -725 488
rect -691 -488 -685 488
rect -731 -500 -685 -488
rect -613 488 -567 500
rect -613 -488 -607 488
rect -573 -488 -567 488
rect -613 -500 -567 -488
rect -495 488 -449 500
rect -495 -488 -489 488
rect -455 -488 -449 488
rect -495 -500 -449 -488
rect -377 488 -331 500
rect -377 -488 -371 488
rect -337 -488 -331 488
rect -377 -500 -331 -488
rect -259 488 -213 500
rect -259 -488 -253 488
rect -219 -488 -213 488
rect -259 -500 -213 -488
rect -141 488 -95 500
rect -141 -488 -135 488
rect -101 -488 -95 488
rect -141 -500 -95 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 95 488 141 500
rect 95 -488 101 488
rect 135 -488 141 488
rect 95 -500 141 -488
rect 213 488 259 500
rect 213 -488 219 488
rect 253 -488 259 488
rect 213 -500 259 -488
rect 331 488 377 500
rect 331 -488 337 488
rect 371 -488 377 488
rect 331 -500 377 -488
rect 449 488 495 500
rect 449 -488 455 488
rect 489 -488 495 488
rect 449 -500 495 -488
rect 567 488 613 500
rect 567 -488 573 488
rect 607 -488 613 488
rect 567 -500 613 -488
rect 685 488 731 500
rect 685 -488 691 488
rect 725 -488 731 488
rect 685 -500 731 -488
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.3 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
