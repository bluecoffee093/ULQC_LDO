** sch_path: /foss/designs/ulqc_ldo/repo/ULQC_LDO/xschem/untitled.sch
**.subckt untitled
x1 IN VSS VSS VDD VDD OUT sky130_fd_sc_hd__clkinv_2
V1 VDD VSS 1.8
.save i(v1)
V2 IN VSS 0
.save i(v2)
V4 VSS GND 0
.save i(v4)
**** begin user architecture code

.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.saveall
.dc temp -40 120



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.saveall
.control
dc V2 0 1.8 0.01
plot v(OUT)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
