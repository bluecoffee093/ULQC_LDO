magic
tech sky130A
magscale 1 2
timestamp 1697815432
<< nmos >>
rect -2035 -500 -1835 500
rect -1777 -500 -1577 500
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
rect 1577 -500 1777 500
rect 1835 -500 2035 500
<< ndiff >>
rect -2093 488 -2035 500
rect -2093 -488 -2081 488
rect -2047 -488 -2035 488
rect -2093 -500 -2035 -488
rect -1835 488 -1777 500
rect -1835 -488 -1823 488
rect -1789 -488 -1777 488
rect -1835 -500 -1777 -488
rect -1577 488 -1519 500
rect -1577 -488 -1565 488
rect -1531 -488 -1519 488
rect -1577 -500 -1519 -488
rect -1319 488 -1261 500
rect -1319 -488 -1307 488
rect -1273 -488 -1261 488
rect -1319 -500 -1261 -488
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
rect 1261 488 1319 500
rect 1261 -488 1273 488
rect 1307 -488 1319 488
rect 1261 -500 1319 -488
rect 1519 488 1577 500
rect 1519 -488 1531 488
rect 1565 -488 1577 488
rect 1519 -500 1577 -488
rect 1777 488 1835 500
rect 1777 -488 1789 488
rect 1823 -488 1835 488
rect 1777 -500 1835 -488
rect 2035 488 2093 500
rect 2035 -488 2047 488
rect 2081 -488 2093 488
rect 2035 -500 2093 -488
<< ndiffc >>
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
<< poly >>
rect -2035 500 -1835 526
rect -1777 500 -1577 526
rect -1519 500 -1319 526
rect -1261 500 -1061 526
rect -1003 500 -803 526
rect -745 500 -545 526
rect -487 500 -287 526
rect -229 500 -29 526
rect 29 500 229 526
rect 287 500 487 526
rect 545 500 745 526
rect 803 500 1003 526
rect 1061 500 1261 526
rect 1319 500 1519 526
rect 1577 500 1777 526
rect 1835 500 2035 526
rect -2035 -526 -1835 -500
rect -1777 -526 -1577 -500
rect -1519 -526 -1319 -500
rect -1261 -526 -1061 -500
rect -1003 -526 -803 -500
rect -745 -526 -545 -500
rect -487 -526 -287 -500
rect -229 -526 -29 -500
rect 29 -526 229 -500
rect 287 -526 487 -500
rect 545 -526 745 -500
rect 803 -526 1003 -500
rect 1061 -526 1261 -500
rect 1319 -526 1519 -500
rect 1577 -526 1777 -500
rect 1835 -526 2035 -500
<< locali >>
rect -2081 488 -2047 504
rect -2081 -504 -2047 -488
rect -1823 488 -1789 504
rect -1823 -504 -1789 -488
rect -1565 488 -1531 504
rect -1565 -504 -1531 -488
rect -1307 488 -1273 504
rect -1307 -504 -1273 -488
rect -1049 488 -1015 504
rect -1049 -504 -1015 -488
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -504 1049 -488
rect 1273 488 1307 504
rect 1273 -504 1307 -488
rect 1531 488 1565 504
rect 1531 -504 1565 -488
rect 1789 488 1823 504
rect 1789 -504 1823 -488
rect 2047 488 2081 504
rect 2047 -504 2081 -488
<< viali >>
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
<< metal1 >>
rect -2087 488 -2041 500
rect -2087 -488 -2081 488
rect -2047 -488 -2041 488
rect -2087 -500 -2041 -488
rect -1829 488 -1783 500
rect -1829 -488 -1823 488
rect -1789 -488 -1783 488
rect -1829 -500 -1783 -488
rect -1571 488 -1525 500
rect -1571 -488 -1565 488
rect -1531 -488 -1525 488
rect -1571 -500 -1525 -488
rect -1313 488 -1267 500
rect -1313 -488 -1307 488
rect -1273 -488 -1267 488
rect -1313 -500 -1267 -488
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect 1267 488 1313 500
rect 1267 -488 1273 488
rect 1307 -488 1313 488
rect 1267 -500 1313 -488
rect 1525 488 1571 500
rect 1525 -488 1531 488
rect 1565 -488 1571 488
rect 1525 -500 1571 -488
rect 1783 488 1829 500
rect 1783 -488 1789 488
rect 1823 -488 1829 488
rect 1783 -500 1829 -488
rect 2041 488 2087 500
rect 2041 -488 2047 488
rect 2081 -488 2087 488
rect 2041 -500 2087 -488
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 1 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
