magic
tech sky130A
magscale 1 2
timestamp 1697926267
<< pwell >>
rect -5457 -3210 5457 3210
<< nmoslvt >>
rect -5261 -3000 -4261 3000
rect -4203 -3000 -3203 3000
rect -3145 -3000 -2145 3000
rect -2087 -3000 -1087 3000
rect -1029 -3000 -29 3000
rect 29 -3000 1029 3000
rect 1087 -3000 2087 3000
rect 2145 -3000 3145 3000
rect 3203 -3000 4203 3000
rect 4261 -3000 5261 3000
<< ndiff >>
rect -5319 2988 -5261 3000
rect -5319 -2988 -5307 2988
rect -5273 -2988 -5261 2988
rect -5319 -3000 -5261 -2988
rect -4261 2988 -4203 3000
rect -4261 -2988 -4249 2988
rect -4215 -2988 -4203 2988
rect -4261 -3000 -4203 -2988
rect -3203 2988 -3145 3000
rect -3203 -2988 -3191 2988
rect -3157 -2988 -3145 2988
rect -3203 -3000 -3145 -2988
rect -2145 2988 -2087 3000
rect -2145 -2988 -2133 2988
rect -2099 -2988 -2087 2988
rect -2145 -3000 -2087 -2988
rect -1087 2988 -1029 3000
rect -1087 -2988 -1075 2988
rect -1041 -2988 -1029 2988
rect -1087 -3000 -1029 -2988
rect -29 2988 29 3000
rect -29 -2988 -17 2988
rect 17 -2988 29 2988
rect -29 -3000 29 -2988
rect 1029 2988 1087 3000
rect 1029 -2988 1041 2988
rect 1075 -2988 1087 2988
rect 1029 -3000 1087 -2988
rect 2087 2988 2145 3000
rect 2087 -2988 2099 2988
rect 2133 -2988 2145 2988
rect 2087 -3000 2145 -2988
rect 3145 2988 3203 3000
rect 3145 -2988 3157 2988
rect 3191 -2988 3203 2988
rect 3145 -3000 3203 -2988
rect 4203 2988 4261 3000
rect 4203 -2988 4215 2988
rect 4249 -2988 4261 2988
rect 4203 -3000 4261 -2988
rect 5261 2988 5319 3000
rect 5261 -2988 5273 2988
rect 5307 -2988 5319 2988
rect 5261 -3000 5319 -2988
<< ndiffc >>
rect -5307 -2988 -5273 2988
rect -4249 -2988 -4215 2988
rect -3191 -2988 -3157 2988
rect -2133 -2988 -2099 2988
rect -1075 -2988 -1041 2988
rect -17 -2988 17 2988
rect 1041 -2988 1075 2988
rect 2099 -2988 2133 2988
rect 3157 -2988 3191 2988
rect 4215 -2988 4249 2988
rect 5273 -2988 5307 2988
<< psubdiff >>
rect -5421 3140 -5325 3174
rect 5325 3140 5421 3174
rect -5421 3078 -5387 3140
rect 5387 3078 5421 3140
rect -5421 -3140 -5387 -3078
rect 5387 -3140 5421 -3078
rect -5421 -3174 -5325 -3140
rect 5325 -3174 5421 -3140
<< psubdiffcont >>
rect -5325 3140 5325 3174
rect -5421 -3078 -5387 3078
rect 5387 -3078 5421 3078
rect -5325 -3174 5325 -3140
<< poly >>
rect -5261 3072 -4261 3088
rect -5261 3038 -5245 3072
rect -4277 3038 -4261 3072
rect -5261 3000 -4261 3038
rect -4203 3072 -3203 3088
rect -4203 3038 -4187 3072
rect -3219 3038 -3203 3072
rect -4203 3000 -3203 3038
rect -3145 3072 -2145 3088
rect -3145 3038 -3129 3072
rect -2161 3038 -2145 3072
rect -3145 3000 -2145 3038
rect -2087 3072 -1087 3088
rect -2087 3038 -2071 3072
rect -1103 3038 -1087 3072
rect -2087 3000 -1087 3038
rect -1029 3072 -29 3088
rect -1029 3038 -1013 3072
rect -45 3038 -29 3072
rect -1029 3000 -29 3038
rect 29 3072 1029 3088
rect 29 3038 45 3072
rect 1013 3038 1029 3072
rect 29 3000 1029 3038
rect 1087 3072 2087 3088
rect 1087 3038 1103 3072
rect 2071 3038 2087 3072
rect 1087 3000 2087 3038
rect 2145 3072 3145 3088
rect 2145 3038 2161 3072
rect 3129 3038 3145 3072
rect 2145 3000 3145 3038
rect 3203 3072 4203 3088
rect 3203 3038 3219 3072
rect 4187 3038 4203 3072
rect 3203 3000 4203 3038
rect 4261 3072 5261 3088
rect 4261 3038 4277 3072
rect 5245 3038 5261 3072
rect 4261 3000 5261 3038
rect -5261 -3038 -4261 -3000
rect -5261 -3072 -5245 -3038
rect -4277 -3072 -4261 -3038
rect -5261 -3088 -4261 -3072
rect -4203 -3038 -3203 -3000
rect -4203 -3072 -4187 -3038
rect -3219 -3072 -3203 -3038
rect -4203 -3088 -3203 -3072
rect -3145 -3038 -2145 -3000
rect -3145 -3072 -3129 -3038
rect -2161 -3072 -2145 -3038
rect -3145 -3088 -2145 -3072
rect -2087 -3038 -1087 -3000
rect -2087 -3072 -2071 -3038
rect -1103 -3072 -1087 -3038
rect -2087 -3088 -1087 -3072
rect -1029 -3038 -29 -3000
rect -1029 -3072 -1013 -3038
rect -45 -3072 -29 -3038
rect -1029 -3088 -29 -3072
rect 29 -3038 1029 -3000
rect 29 -3072 45 -3038
rect 1013 -3072 1029 -3038
rect 29 -3088 1029 -3072
rect 1087 -3038 2087 -3000
rect 1087 -3072 1103 -3038
rect 2071 -3072 2087 -3038
rect 1087 -3088 2087 -3072
rect 2145 -3038 3145 -3000
rect 2145 -3072 2161 -3038
rect 3129 -3072 3145 -3038
rect 2145 -3088 3145 -3072
rect 3203 -3038 4203 -3000
rect 3203 -3072 3219 -3038
rect 4187 -3072 4203 -3038
rect 3203 -3088 4203 -3072
rect 4261 -3038 5261 -3000
rect 4261 -3072 4277 -3038
rect 5245 -3072 5261 -3038
rect 4261 -3088 5261 -3072
<< polycont >>
rect -5245 3038 -4277 3072
rect -4187 3038 -3219 3072
rect -3129 3038 -2161 3072
rect -2071 3038 -1103 3072
rect -1013 3038 -45 3072
rect 45 3038 1013 3072
rect 1103 3038 2071 3072
rect 2161 3038 3129 3072
rect 3219 3038 4187 3072
rect 4277 3038 5245 3072
rect -5245 -3072 -4277 -3038
rect -4187 -3072 -3219 -3038
rect -3129 -3072 -2161 -3038
rect -2071 -3072 -1103 -3038
rect -1013 -3072 -45 -3038
rect 45 -3072 1013 -3038
rect 1103 -3072 2071 -3038
rect 2161 -3072 3129 -3038
rect 3219 -3072 4187 -3038
rect 4277 -3072 5245 -3038
<< locali >>
rect -5421 3140 -5325 3174
rect 5325 3140 5421 3174
rect -5421 3078 -5387 3140
rect 5387 3078 5421 3140
rect -5261 3038 -5245 3072
rect -4277 3038 -4261 3072
rect -4203 3038 -4187 3072
rect -3219 3038 -3203 3072
rect -3145 3038 -3129 3072
rect -2161 3038 -2145 3072
rect -2087 3038 -2071 3072
rect -1103 3038 -1087 3072
rect -1029 3038 -1013 3072
rect -45 3038 -29 3072
rect 29 3038 45 3072
rect 1013 3038 1029 3072
rect 1087 3038 1103 3072
rect 2071 3038 2087 3072
rect 2145 3038 2161 3072
rect 3129 3038 3145 3072
rect 3203 3038 3219 3072
rect 4187 3038 4203 3072
rect 4261 3038 4277 3072
rect 5245 3038 5261 3072
rect -5307 2988 -5273 3004
rect -5307 -3004 -5273 -2988
rect -4249 2988 -4215 3004
rect -4249 -3004 -4215 -2988
rect -3191 2988 -3157 3004
rect -3191 -3004 -3157 -2988
rect -2133 2988 -2099 3004
rect -2133 -3004 -2099 -2988
rect -1075 2988 -1041 3004
rect -1075 -3004 -1041 -2988
rect -17 2988 17 3004
rect -17 -3004 17 -2988
rect 1041 2988 1075 3004
rect 1041 -3004 1075 -2988
rect 2099 2988 2133 3004
rect 2099 -3004 2133 -2988
rect 3157 2988 3191 3004
rect 3157 -3004 3191 -2988
rect 4215 2988 4249 3004
rect 4215 -3004 4249 -2988
rect 5273 2988 5307 3004
rect 5273 -3004 5307 -2988
rect -5261 -3072 -5245 -3038
rect -4277 -3072 -4261 -3038
rect -4203 -3072 -4187 -3038
rect -3219 -3072 -3203 -3038
rect -3145 -3072 -3129 -3038
rect -2161 -3072 -2145 -3038
rect -2087 -3072 -2071 -3038
rect -1103 -3072 -1087 -3038
rect -1029 -3072 -1013 -3038
rect -45 -3072 -29 -3038
rect 29 -3072 45 -3038
rect 1013 -3072 1029 -3038
rect 1087 -3072 1103 -3038
rect 2071 -3072 2087 -3038
rect 2145 -3072 2161 -3038
rect 3129 -3072 3145 -3038
rect 3203 -3072 3219 -3038
rect 4187 -3072 4203 -3038
rect 4261 -3072 4277 -3038
rect 5245 -3072 5261 -3038
rect -5421 -3140 -5387 -3078
rect 5387 -3140 5421 -3078
rect -5421 -3174 -5325 -3140
rect 5325 -3174 5421 -3140
<< viali >>
rect -5245 3038 -4277 3072
rect -4187 3038 -3219 3072
rect -3129 3038 -2161 3072
rect -2071 3038 -1103 3072
rect -1013 3038 -45 3072
rect 45 3038 1013 3072
rect 1103 3038 2071 3072
rect 2161 3038 3129 3072
rect 3219 3038 4187 3072
rect 4277 3038 5245 3072
rect -5307 -2988 -5273 2988
rect -4249 -2988 -4215 2988
rect -3191 -2988 -3157 2988
rect -2133 -2988 -2099 2988
rect -1075 -2988 -1041 2988
rect -17 -2988 17 2988
rect 1041 -2988 1075 2988
rect 2099 -2988 2133 2988
rect 3157 -2988 3191 2988
rect 4215 -2988 4249 2988
rect 5273 -2988 5307 2988
rect -5245 -3072 -4277 -3038
rect -4187 -3072 -3219 -3038
rect -3129 -3072 -2161 -3038
rect -2071 -3072 -1103 -3038
rect -1013 -3072 -45 -3038
rect 45 -3072 1013 -3038
rect 1103 -3072 2071 -3038
rect 2161 -3072 3129 -3038
rect 3219 -3072 4187 -3038
rect 4277 -3072 5245 -3038
<< metal1 >>
rect -5257 3072 -4265 3078
rect -5257 3038 -5245 3072
rect -4277 3038 -4265 3072
rect -5257 3032 -4265 3038
rect -4199 3072 -3207 3078
rect -4199 3038 -4187 3072
rect -3219 3038 -3207 3072
rect -4199 3032 -3207 3038
rect -3141 3072 -2149 3078
rect -3141 3038 -3129 3072
rect -2161 3038 -2149 3072
rect -3141 3032 -2149 3038
rect -2083 3072 -1091 3078
rect -2083 3038 -2071 3072
rect -1103 3038 -1091 3072
rect -2083 3032 -1091 3038
rect -1025 3072 -33 3078
rect -1025 3038 -1013 3072
rect -45 3038 -33 3072
rect -1025 3032 -33 3038
rect 33 3072 1025 3078
rect 33 3038 45 3072
rect 1013 3038 1025 3072
rect 33 3032 1025 3038
rect 1091 3072 2083 3078
rect 1091 3038 1103 3072
rect 2071 3038 2083 3072
rect 1091 3032 2083 3038
rect 2149 3072 3141 3078
rect 2149 3038 2161 3072
rect 3129 3038 3141 3072
rect 2149 3032 3141 3038
rect 3207 3072 4199 3078
rect 3207 3038 3219 3072
rect 4187 3038 4199 3072
rect 3207 3032 4199 3038
rect 4265 3072 5257 3078
rect 4265 3038 4277 3072
rect 5245 3038 5257 3072
rect 4265 3032 5257 3038
rect -5313 2988 -5267 3000
rect -5313 -2988 -5307 2988
rect -5273 -2988 -5267 2988
rect -5313 -3000 -5267 -2988
rect -4255 2988 -4209 3000
rect -4255 -2988 -4249 2988
rect -4215 -2988 -4209 2988
rect -4255 -3000 -4209 -2988
rect -3197 2988 -3151 3000
rect -3197 -2988 -3191 2988
rect -3157 -2988 -3151 2988
rect -3197 -3000 -3151 -2988
rect -2139 2988 -2093 3000
rect -2139 -2988 -2133 2988
rect -2099 -2988 -2093 2988
rect -2139 -3000 -2093 -2988
rect -1081 2988 -1035 3000
rect -1081 -2988 -1075 2988
rect -1041 -2988 -1035 2988
rect -1081 -3000 -1035 -2988
rect -23 2988 23 3000
rect -23 -2988 -17 2988
rect 17 -2988 23 2988
rect -23 -3000 23 -2988
rect 1035 2988 1081 3000
rect 1035 -2988 1041 2988
rect 1075 -2988 1081 2988
rect 1035 -3000 1081 -2988
rect 2093 2988 2139 3000
rect 2093 -2988 2099 2988
rect 2133 -2988 2139 2988
rect 2093 -3000 2139 -2988
rect 3151 2988 3197 3000
rect 3151 -2988 3157 2988
rect 3191 -2988 3197 2988
rect 3151 -3000 3197 -2988
rect 4209 2988 4255 3000
rect 4209 -2988 4215 2988
rect 4249 -2988 4255 2988
rect 4209 -3000 4255 -2988
rect 5267 2988 5313 3000
rect 5267 -2988 5273 2988
rect 5307 -2988 5313 2988
rect 5267 -3000 5313 -2988
rect -5257 -3038 -4265 -3032
rect -5257 -3072 -5245 -3038
rect -4277 -3072 -4265 -3038
rect -5257 -3078 -4265 -3072
rect -4199 -3038 -3207 -3032
rect -4199 -3072 -4187 -3038
rect -3219 -3072 -3207 -3038
rect -4199 -3078 -3207 -3072
rect -3141 -3038 -2149 -3032
rect -3141 -3072 -3129 -3038
rect -2161 -3072 -2149 -3038
rect -3141 -3078 -2149 -3072
rect -2083 -3038 -1091 -3032
rect -2083 -3072 -2071 -3038
rect -1103 -3072 -1091 -3038
rect -2083 -3078 -1091 -3072
rect -1025 -3038 -33 -3032
rect -1025 -3072 -1013 -3038
rect -45 -3072 -33 -3038
rect -1025 -3078 -33 -3072
rect 33 -3038 1025 -3032
rect 33 -3072 45 -3038
rect 1013 -3072 1025 -3038
rect 33 -3078 1025 -3072
rect 1091 -3038 2083 -3032
rect 1091 -3072 1103 -3038
rect 2071 -3072 2083 -3038
rect 1091 -3078 2083 -3072
rect 2149 -3038 3141 -3032
rect 2149 -3072 2161 -3038
rect 3129 -3072 3141 -3038
rect 2149 -3078 3141 -3072
rect 3207 -3038 4199 -3032
rect 3207 -3072 3219 -3038
rect 4187 -3072 4199 -3038
rect 3207 -3078 4199 -3072
rect 4265 -3038 5257 -3032
rect 4265 -3072 4277 -3038
rect 5245 -3072 5257 -3038
rect 4265 -3078 5257 -3072
<< properties >>
string FIXED_BBOX -5404 -3157 5404 3157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 30.0 l 5.0 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
