** sch_path: /foss/designs/ulqc_ldo/repo/ULQC_LDO/xschem/bandgap.sch
.subckt bandgap BGR_OUT VDD VSS BGRT1 BGRT2
*.PININFO BGR_OUT:O VDD:I VSS:I BGRT1:I BGRT2:I
XM7 net1 net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=60 nf=1 m=8
XM8 net2 net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=60 nf=1 m=8
XM9 net2 net1 v2 VSS sky130_fd_pr__nfet_01v8_lvt L=10 W=60 nf=1 m=8
XM10 net1 net1 v1 VSS sky130_fd_pr__nfet_01v8_lvt L=10 W=60 nf=1 m=8
XQ4 VSS VSS net3 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=8
XQ5 VSS VSS v1 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
XM11 BGR_OUT net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=60 nf=1 m=8
x9 VSS_60 VCC_60 VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x15 VSS_70 VCC_70 VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x17 VSS_80 VCC_80 VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x18 VSS_85 VCC_85 VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x19 net5 BGRT1 VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x20 net4 BGRT2 VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
XR7 net11 BGR_OUT VSS sky130_fd_pr__res_high_po_0p35 L=15 mult=1 m=1
XM12 net2 net2 net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=10 nf=1 m=1
XR8 net3 v2 VSS sky130_fd_pr__res_high_po_0p35 L=8.8 mult=1 m=1
XR9 net6 net7 VSS sky130_fd_pr__res_high_po_0p35 L=19 mult=1 m=1
x22 VDD BGRT1 VCC_60 BGRT2 VSS and_gate
x23 VDD net5 VCC_70 net4 VSS and_gate
x24 VDD net5 VCC_80 BGRT2 VSS and_gate
x25 VDD BGRT1 VCC_85 net4 VSS and_gate
XR10 net8 net6 VSS sky130_fd_pr__res_high_po_0p35 L=22 mult=1 m=1
XR11 net9 net8 VSS sky130_fd_pr__res_high_po_0p35 L=25.3 mult=1 m=1
XR12 net10 net9 VSS sky130_fd_pr__res_high_po_0p35 L=27 mult=1 m=1
XQ6 VSS VSS net10 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
x1 net6 net7 VCC_60 VSS_60 VCC VSS passgate_nlvt W_N=1 L_N=0.35 W_P=1 L_P=0.35 m=1
x2 net8 net6 VCC_70 VSS_70 VCC VSS passgate_nlvt W_N=1 L_N=0.35 W_P=1 L_P=0.35 m=1
x3 net9 net8 VCC_80 VSS_80 VCC VSS passgate_nlvt W_N=1 L_N=0.35 W_P=1 L_P=0.35 m=1
x4 net10 net9 VCC_85 VSS_85 VCC VSS passgate_nlvt W_N=1 L_N=0.35 W_P=1 L_P=0.35 m=1
XR1 net12 net11 VSS sky130_fd_pr__res_high_po_0p35 L=15 mult=1 m=1
XR2 net7 net12 VSS sky130_fd_pr__res_high_po_0p35 L=15 mult=1 m=1
.ends

* expanding   symbol:  sky130_tests/not.sym # of pins=2
** sym_path: /foss/pdks/sky130A/libs.tech/xschem/sky130_tests/not.sym
** sch_path: /foss/pdks/sky130A/libs.tech/xschem/sky130_tests/not.sch
.subckt not y a VCCPIN VSSPIN     W_N=1 L_N=0.15 W_P=2 L_P=0.15
*.PININFO y:O a:I
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 m=1
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 m=1
.ends


* expanding   symbol:  /foss/designs/ulqc_ldo/repo/ULQC_LDO/xschem/and_gate.sym # of pins=5
** sym_path: /foss/designs/ulqc_ldo/repo/ULQC_LDO/xschem/and_gate.sym
** sch_path: /foss/designs/ulqc_ldo/repo/ULQC_LDO/xschem/and_gate.sch
.subckt and_gate VDD A OUT B VSS
*.PININFO OUT:O A:I B:I VDD:I VSS:I
XM1 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 net1 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 net1 A net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net2 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 OUT net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  sky130_tests/passgate_nlvt.sym # of pins=4
** sym_path: /foss/pdks/sky130A/libs.tech/xschem/sky130_tests/passgate_nlvt.sym
** sch_path: /foss/pdks/sky130A/libs.tech/xschem/sky130_tests/passgate_nlvt.sch
.subckt passgate_nlvt Z A GP GN VCCBPIN VSSBPIN  W_N=1 L_N=0.35 W_P=1 L_P=0.35
*.PININFO A:B Z:B GP:I GN:I
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8_lvt L=L_N W=W_N nf=1 m=1
XM2 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8_lvt L=L_P W=W_P nf=1 m=1
* noconn VCCBPIN
* noconn VSSBPIN
.ends

.end
