magic
tech sky130A
magscale 1 2
timestamp 1697796765
<< error_p >>
rect -2765 3290 -2707 3296
rect -2573 3290 -2515 3296
rect -2381 3290 -2323 3296
rect -2189 3290 -2131 3296
rect -1997 3290 -1939 3296
rect -1805 3290 -1747 3296
rect -1613 3290 -1555 3296
rect -1421 3290 -1363 3296
rect -1229 3290 -1171 3296
rect -1037 3290 -979 3296
rect -845 3290 -787 3296
rect -653 3290 -595 3296
rect -461 3290 -403 3296
rect -269 3290 -211 3296
rect -77 3290 -19 3296
rect 115 3290 173 3296
rect 307 3290 365 3296
rect 499 3290 557 3296
rect 691 3290 749 3296
rect 883 3290 941 3296
rect 1075 3290 1133 3296
rect 1267 3290 1325 3296
rect 1459 3290 1517 3296
rect 1651 3290 1709 3296
rect 1843 3290 1901 3296
rect 2035 3290 2093 3296
rect 2227 3290 2285 3296
rect 2419 3290 2477 3296
rect 2611 3290 2669 3296
rect 2803 3290 2861 3296
rect -2765 3256 -2753 3290
rect -2573 3256 -2561 3290
rect -2381 3256 -2369 3290
rect -2189 3256 -2177 3290
rect -1997 3256 -1985 3290
rect -1805 3256 -1793 3290
rect -1613 3256 -1601 3290
rect -1421 3256 -1409 3290
rect -1229 3256 -1217 3290
rect -1037 3256 -1025 3290
rect -845 3256 -833 3290
rect -653 3256 -641 3290
rect -461 3256 -449 3290
rect -269 3256 -257 3290
rect -77 3256 -65 3290
rect 115 3256 127 3290
rect 307 3256 319 3290
rect 499 3256 511 3290
rect 691 3256 703 3290
rect 883 3256 895 3290
rect 1075 3256 1087 3290
rect 1267 3256 1279 3290
rect 1459 3256 1471 3290
rect 1651 3256 1663 3290
rect 1843 3256 1855 3290
rect 2035 3256 2047 3290
rect 2227 3256 2239 3290
rect 2419 3256 2431 3290
rect 2611 3256 2623 3290
rect 2803 3256 2815 3290
rect -2765 3250 -2707 3256
rect -2573 3250 -2515 3256
rect -2381 3250 -2323 3256
rect -2189 3250 -2131 3256
rect -1997 3250 -1939 3256
rect -1805 3250 -1747 3256
rect -1613 3250 -1555 3256
rect -1421 3250 -1363 3256
rect -1229 3250 -1171 3256
rect -1037 3250 -979 3256
rect -845 3250 -787 3256
rect -653 3250 -595 3256
rect -461 3250 -403 3256
rect -269 3250 -211 3256
rect -77 3250 -19 3256
rect 115 3250 173 3256
rect 307 3250 365 3256
rect 499 3250 557 3256
rect 691 3250 749 3256
rect 883 3250 941 3256
rect 1075 3250 1133 3256
rect 1267 3250 1325 3256
rect 1459 3250 1517 3256
rect 1651 3250 1709 3256
rect 1843 3250 1901 3256
rect 2035 3250 2093 3256
rect 2227 3250 2285 3256
rect 2419 3250 2477 3256
rect 2611 3250 2669 3256
rect 2803 3250 2861 3256
rect -2861 1180 -2803 1186
rect -2669 1180 -2611 1186
rect -2477 1180 -2419 1186
rect -2285 1180 -2227 1186
rect -2093 1180 -2035 1186
rect -1901 1180 -1843 1186
rect -1709 1180 -1651 1186
rect -1517 1180 -1459 1186
rect -1325 1180 -1267 1186
rect -1133 1180 -1075 1186
rect -941 1180 -883 1186
rect -749 1180 -691 1186
rect -557 1180 -499 1186
rect -365 1180 -307 1186
rect -173 1180 -115 1186
rect 19 1180 77 1186
rect 211 1180 269 1186
rect 403 1180 461 1186
rect 595 1180 653 1186
rect 787 1180 845 1186
rect 979 1180 1037 1186
rect 1171 1180 1229 1186
rect 1363 1180 1421 1186
rect 1555 1180 1613 1186
rect 1747 1180 1805 1186
rect 1939 1180 1997 1186
rect 2131 1180 2189 1186
rect 2323 1180 2381 1186
rect 2515 1180 2573 1186
rect 2707 1180 2765 1186
rect -2861 1146 -2849 1180
rect -2669 1146 -2657 1180
rect -2477 1146 -2465 1180
rect -2285 1146 -2273 1180
rect -2093 1146 -2081 1180
rect -1901 1146 -1889 1180
rect -1709 1146 -1697 1180
rect -1517 1146 -1505 1180
rect -1325 1146 -1313 1180
rect -1133 1146 -1121 1180
rect -941 1146 -929 1180
rect -749 1146 -737 1180
rect -557 1146 -545 1180
rect -365 1146 -353 1180
rect -173 1146 -161 1180
rect 19 1146 31 1180
rect 211 1146 223 1180
rect 403 1146 415 1180
rect 595 1146 607 1180
rect 787 1146 799 1180
rect 979 1146 991 1180
rect 1171 1146 1183 1180
rect 1363 1146 1375 1180
rect 1555 1146 1567 1180
rect 1747 1146 1759 1180
rect 1939 1146 1951 1180
rect 2131 1146 2143 1180
rect 2323 1146 2335 1180
rect 2515 1146 2527 1180
rect 2707 1146 2719 1180
rect -2861 1140 -2803 1146
rect -2669 1140 -2611 1146
rect -2477 1140 -2419 1146
rect -2285 1140 -2227 1146
rect -2093 1140 -2035 1146
rect -1901 1140 -1843 1146
rect -1709 1140 -1651 1146
rect -1517 1140 -1459 1146
rect -1325 1140 -1267 1146
rect -1133 1140 -1075 1146
rect -941 1140 -883 1146
rect -749 1140 -691 1146
rect -557 1140 -499 1146
rect -365 1140 -307 1146
rect -173 1140 -115 1146
rect 19 1140 77 1146
rect 211 1140 269 1146
rect 403 1140 461 1146
rect 595 1140 653 1146
rect 787 1140 845 1146
rect 979 1140 1037 1146
rect 1171 1140 1229 1146
rect 1363 1140 1421 1146
rect 1555 1140 1613 1146
rect 1747 1140 1805 1146
rect 1939 1140 1997 1146
rect 2131 1140 2189 1146
rect 2323 1140 2381 1146
rect 2515 1140 2573 1146
rect 2707 1140 2765 1146
rect -2861 1072 -2803 1078
rect -2669 1072 -2611 1078
rect -2477 1072 -2419 1078
rect -2285 1072 -2227 1078
rect -2093 1072 -2035 1078
rect -1901 1072 -1843 1078
rect -1709 1072 -1651 1078
rect -1517 1072 -1459 1078
rect -1325 1072 -1267 1078
rect -1133 1072 -1075 1078
rect -941 1072 -883 1078
rect -749 1072 -691 1078
rect -557 1072 -499 1078
rect -365 1072 -307 1078
rect -173 1072 -115 1078
rect 19 1072 77 1078
rect 211 1072 269 1078
rect 403 1072 461 1078
rect 595 1072 653 1078
rect 787 1072 845 1078
rect 979 1072 1037 1078
rect 1171 1072 1229 1078
rect 1363 1072 1421 1078
rect 1555 1072 1613 1078
rect 1747 1072 1805 1078
rect 1939 1072 1997 1078
rect 2131 1072 2189 1078
rect 2323 1072 2381 1078
rect 2515 1072 2573 1078
rect 2707 1072 2765 1078
rect -2861 1038 -2849 1072
rect -2669 1038 -2657 1072
rect -2477 1038 -2465 1072
rect -2285 1038 -2273 1072
rect -2093 1038 -2081 1072
rect -1901 1038 -1889 1072
rect -1709 1038 -1697 1072
rect -1517 1038 -1505 1072
rect -1325 1038 -1313 1072
rect -1133 1038 -1121 1072
rect -941 1038 -929 1072
rect -749 1038 -737 1072
rect -557 1038 -545 1072
rect -365 1038 -353 1072
rect -173 1038 -161 1072
rect 19 1038 31 1072
rect 211 1038 223 1072
rect 403 1038 415 1072
rect 595 1038 607 1072
rect 787 1038 799 1072
rect 979 1038 991 1072
rect 1171 1038 1183 1072
rect 1363 1038 1375 1072
rect 1555 1038 1567 1072
rect 1747 1038 1759 1072
rect 1939 1038 1951 1072
rect 2131 1038 2143 1072
rect 2323 1038 2335 1072
rect 2515 1038 2527 1072
rect 2707 1038 2719 1072
rect -2861 1032 -2803 1038
rect -2669 1032 -2611 1038
rect -2477 1032 -2419 1038
rect -2285 1032 -2227 1038
rect -2093 1032 -2035 1038
rect -1901 1032 -1843 1038
rect -1709 1032 -1651 1038
rect -1517 1032 -1459 1038
rect -1325 1032 -1267 1038
rect -1133 1032 -1075 1038
rect -941 1032 -883 1038
rect -749 1032 -691 1038
rect -557 1032 -499 1038
rect -365 1032 -307 1038
rect -173 1032 -115 1038
rect 19 1032 77 1038
rect 211 1032 269 1038
rect 403 1032 461 1038
rect 595 1032 653 1038
rect 787 1032 845 1038
rect 979 1032 1037 1038
rect 1171 1032 1229 1038
rect 1363 1032 1421 1038
rect 1555 1032 1613 1038
rect 1747 1032 1805 1038
rect 1939 1032 1997 1038
rect 2131 1032 2189 1038
rect 2323 1032 2381 1038
rect 2515 1032 2573 1038
rect 2707 1032 2765 1038
rect -2765 -1038 -2707 -1032
rect -2573 -1038 -2515 -1032
rect -2381 -1038 -2323 -1032
rect -2189 -1038 -2131 -1032
rect -1997 -1038 -1939 -1032
rect -1805 -1038 -1747 -1032
rect -1613 -1038 -1555 -1032
rect -1421 -1038 -1363 -1032
rect -1229 -1038 -1171 -1032
rect -1037 -1038 -979 -1032
rect -845 -1038 -787 -1032
rect -653 -1038 -595 -1032
rect -461 -1038 -403 -1032
rect -269 -1038 -211 -1032
rect -77 -1038 -19 -1032
rect 115 -1038 173 -1032
rect 307 -1038 365 -1032
rect 499 -1038 557 -1032
rect 691 -1038 749 -1032
rect 883 -1038 941 -1032
rect 1075 -1038 1133 -1032
rect 1267 -1038 1325 -1032
rect 1459 -1038 1517 -1032
rect 1651 -1038 1709 -1032
rect 1843 -1038 1901 -1032
rect 2035 -1038 2093 -1032
rect 2227 -1038 2285 -1032
rect 2419 -1038 2477 -1032
rect 2611 -1038 2669 -1032
rect 2803 -1038 2861 -1032
rect -2765 -1072 -2753 -1038
rect -2573 -1072 -2561 -1038
rect -2381 -1072 -2369 -1038
rect -2189 -1072 -2177 -1038
rect -1997 -1072 -1985 -1038
rect -1805 -1072 -1793 -1038
rect -1613 -1072 -1601 -1038
rect -1421 -1072 -1409 -1038
rect -1229 -1072 -1217 -1038
rect -1037 -1072 -1025 -1038
rect -845 -1072 -833 -1038
rect -653 -1072 -641 -1038
rect -461 -1072 -449 -1038
rect -269 -1072 -257 -1038
rect -77 -1072 -65 -1038
rect 115 -1072 127 -1038
rect 307 -1072 319 -1038
rect 499 -1072 511 -1038
rect 691 -1072 703 -1038
rect 883 -1072 895 -1038
rect 1075 -1072 1087 -1038
rect 1267 -1072 1279 -1038
rect 1459 -1072 1471 -1038
rect 1651 -1072 1663 -1038
rect 1843 -1072 1855 -1038
rect 2035 -1072 2047 -1038
rect 2227 -1072 2239 -1038
rect 2419 -1072 2431 -1038
rect 2611 -1072 2623 -1038
rect 2803 -1072 2815 -1038
rect -2765 -1078 -2707 -1072
rect -2573 -1078 -2515 -1072
rect -2381 -1078 -2323 -1072
rect -2189 -1078 -2131 -1072
rect -1997 -1078 -1939 -1072
rect -1805 -1078 -1747 -1072
rect -1613 -1078 -1555 -1072
rect -1421 -1078 -1363 -1072
rect -1229 -1078 -1171 -1072
rect -1037 -1078 -979 -1072
rect -845 -1078 -787 -1072
rect -653 -1078 -595 -1072
rect -461 -1078 -403 -1072
rect -269 -1078 -211 -1072
rect -77 -1078 -19 -1072
rect 115 -1078 173 -1072
rect 307 -1078 365 -1072
rect 499 -1078 557 -1072
rect 691 -1078 749 -1072
rect 883 -1078 941 -1072
rect 1075 -1078 1133 -1072
rect 1267 -1078 1325 -1072
rect 1459 -1078 1517 -1072
rect 1651 -1078 1709 -1072
rect 1843 -1078 1901 -1072
rect 2035 -1078 2093 -1072
rect 2227 -1078 2285 -1072
rect 2419 -1078 2477 -1072
rect 2611 -1078 2669 -1072
rect 2803 -1078 2861 -1072
rect -2765 -1146 -2707 -1140
rect -2573 -1146 -2515 -1140
rect -2381 -1146 -2323 -1140
rect -2189 -1146 -2131 -1140
rect -1997 -1146 -1939 -1140
rect -1805 -1146 -1747 -1140
rect -1613 -1146 -1555 -1140
rect -1421 -1146 -1363 -1140
rect -1229 -1146 -1171 -1140
rect -1037 -1146 -979 -1140
rect -845 -1146 -787 -1140
rect -653 -1146 -595 -1140
rect -461 -1146 -403 -1140
rect -269 -1146 -211 -1140
rect -77 -1146 -19 -1140
rect 115 -1146 173 -1140
rect 307 -1146 365 -1140
rect 499 -1146 557 -1140
rect 691 -1146 749 -1140
rect 883 -1146 941 -1140
rect 1075 -1146 1133 -1140
rect 1267 -1146 1325 -1140
rect 1459 -1146 1517 -1140
rect 1651 -1146 1709 -1140
rect 1843 -1146 1901 -1140
rect 2035 -1146 2093 -1140
rect 2227 -1146 2285 -1140
rect 2419 -1146 2477 -1140
rect 2611 -1146 2669 -1140
rect 2803 -1146 2861 -1140
rect -2765 -1180 -2753 -1146
rect -2573 -1180 -2561 -1146
rect -2381 -1180 -2369 -1146
rect -2189 -1180 -2177 -1146
rect -1997 -1180 -1985 -1146
rect -1805 -1180 -1793 -1146
rect -1613 -1180 -1601 -1146
rect -1421 -1180 -1409 -1146
rect -1229 -1180 -1217 -1146
rect -1037 -1180 -1025 -1146
rect -845 -1180 -833 -1146
rect -653 -1180 -641 -1146
rect -461 -1180 -449 -1146
rect -269 -1180 -257 -1146
rect -77 -1180 -65 -1146
rect 115 -1180 127 -1146
rect 307 -1180 319 -1146
rect 499 -1180 511 -1146
rect 691 -1180 703 -1146
rect 883 -1180 895 -1146
rect 1075 -1180 1087 -1146
rect 1267 -1180 1279 -1146
rect 1459 -1180 1471 -1146
rect 1651 -1180 1663 -1146
rect 1843 -1180 1855 -1146
rect 2035 -1180 2047 -1146
rect 2227 -1180 2239 -1146
rect 2419 -1180 2431 -1146
rect 2611 -1180 2623 -1146
rect 2803 -1180 2815 -1146
rect -2765 -1186 -2707 -1180
rect -2573 -1186 -2515 -1180
rect -2381 -1186 -2323 -1180
rect -2189 -1186 -2131 -1180
rect -1997 -1186 -1939 -1180
rect -1805 -1186 -1747 -1180
rect -1613 -1186 -1555 -1180
rect -1421 -1186 -1363 -1180
rect -1229 -1186 -1171 -1180
rect -1037 -1186 -979 -1180
rect -845 -1186 -787 -1180
rect -653 -1186 -595 -1180
rect -461 -1186 -403 -1180
rect -269 -1186 -211 -1180
rect -77 -1186 -19 -1180
rect 115 -1186 173 -1180
rect 307 -1186 365 -1180
rect 499 -1186 557 -1180
rect 691 -1186 749 -1180
rect 883 -1186 941 -1180
rect 1075 -1186 1133 -1180
rect 1267 -1186 1325 -1180
rect 1459 -1186 1517 -1180
rect 1651 -1186 1709 -1180
rect 1843 -1186 1901 -1180
rect 2035 -1186 2093 -1180
rect 2227 -1186 2285 -1180
rect 2419 -1186 2477 -1180
rect 2611 -1186 2669 -1180
rect 2803 -1186 2861 -1180
rect -2861 -3256 -2803 -3250
rect -2669 -3256 -2611 -3250
rect -2477 -3256 -2419 -3250
rect -2285 -3256 -2227 -3250
rect -2093 -3256 -2035 -3250
rect -1901 -3256 -1843 -3250
rect -1709 -3256 -1651 -3250
rect -1517 -3256 -1459 -3250
rect -1325 -3256 -1267 -3250
rect -1133 -3256 -1075 -3250
rect -941 -3256 -883 -3250
rect -749 -3256 -691 -3250
rect -557 -3256 -499 -3250
rect -365 -3256 -307 -3250
rect -173 -3256 -115 -3250
rect 19 -3256 77 -3250
rect 211 -3256 269 -3250
rect 403 -3256 461 -3250
rect 595 -3256 653 -3250
rect 787 -3256 845 -3250
rect 979 -3256 1037 -3250
rect 1171 -3256 1229 -3250
rect 1363 -3256 1421 -3250
rect 1555 -3256 1613 -3250
rect 1747 -3256 1805 -3250
rect 1939 -3256 1997 -3250
rect 2131 -3256 2189 -3250
rect 2323 -3256 2381 -3250
rect 2515 -3256 2573 -3250
rect 2707 -3256 2765 -3250
rect -2861 -3290 -2849 -3256
rect -2669 -3290 -2657 -3256
rect -2477 -3290 -2465 -3256
rect -2285 -3290 -2273 -3256
rect -2093 -3290 -2081 -3256
rect -1901 -3290 -1889 -3256
rect -1709 -3290 -1697 -3256
rect -1517 -3290 -1505 -3256
rect -1325 -3290 -1313 -3256
rect -1133 -3290 -1121 -3256
rect -941 -3290 -929 -3256
rect -749 -3290 -737 -3256
rect -557 -3290 -545 -3256
rect -365 -3290 -353 -3256
rect -173 -3290 -161 -3256
rect 19 -3290 31 -3256
rect 211 -3290 223 -3256
rect 403 -3290 415 -3256
rect 595 -3290 607 -3256
rect 787 -3290 799 -3256
rect 979 -3290 991 -3256
rect 1171 -3290 1183 -3256
rect 1363 -3290 1375 -3256
rect 1555 -3290 1567 -3256
rect 1747 -3290 1759 -3256
rect 1939 -3290 1951 -3256
rect 2131 -3290 2143 -3256
rect 2323 -3290 2335 -3256
rect 2515 -3290 2527 -3256
rect 2707 -3290 2719 -3256
rect -2861 -3296 -2803 -3290
rect -2669 -3296 -2611 -3290
rect -2477 -3296 -2419 -3290
rect -2285 -3296 -2227 -3290
rect -2093 -3296 -2035 -3290
rect -1901 -3296 -1843 -3290
rect -1709 -3296 -1651 -3290
rect -1517 -3296 -1459 -3290
rect -1325 -3296 -1267 -3290
rect -1133 -3296 -1075 -3290
rect -941 -3296 -883 -3290
rect -749 -3296 -691 -3290
rect -557 -3296 -499 -3290
rect -365 -3296 -307 -3290
rect -173 -3296 -115 -3290
rect 19 -3296 77 -3290
rect 211 -3296 269 -3290
rect 403 -3296 461 -3290
rect 595 -3296 653 -3290
rect 787 -3296 845 -3290
rect 979 -3296 1037 -3290
rect 1171 -3296 1229 -3290
rect 1363 -3296 1421 -3290
rect 1555 -3296 1613 -3290
rect 1747 -3296 1805 -3290
rect 1939 -3296 1997 -3290
rect 2131 -3296 2189 -3290
rect 2323 -3296 2381 -3290
rect 2515 -3296 2573 -3290
rect 2707 -3296 2765 -3290
<< nmoslvt >>
rect -2847 1218 -2817 3218
rect -2751 1218 -2721 3218
rect -2655 1218 -2625 3218
rect -2559 1218 -2529 3218
rect -2463 1218 -2433 3218
rect -2367 1218 -2337 3218
rect -2271 1218 -2241 3218
rect -2175 1218 -2145 3218
rect -2079 1218 -2049 3218
rect -1983 1218 -1953 3218
rect -1887 1218 -1857 3218
rect -1791 1218 -1761 3218
rect -1695 1218 -1665 3218
rect -1599 1218 -1569 3218
rect -1503 1218 -1473 3218
rect -1407 1218 -1377 3218
rect -1311 1218 -1281 3218
rect -1215 1218 -1185 3218
rect -1119 1218 -1089 3218
rect -1023 1218 -993 3218
rect -927 1218 -897 3218
rect -831 1218 -801 3218
rect -735 1218 -705 3218
rect -639 1218 -609 3218
rect -543 1218 -513 3218
rect -447 1218 -417 3218
rect -351 1218 -321 3218
rect -255 1218 -225 3218
rect -159 1218 -129 3218
rect -63 1218 -33 3218
rect 33 1218 63 3218
rect 129 1218 159 3218
rect 225 1218 255 3218
rect 321 1218 351 3218
rect 417 1218 447 3218
rect 513 1218 543 3218
rect 609 1218 639 3218
rect 705 1218 735 3218
rect 801 1218 831 3218
rect 897 1218 927 3218
rect 993 1218 1023 3218
rect 1089 1218 1119 3218
rect 1185 1218 1215 3218
rect 1281 1218 1311 3218
rect 1377 1218 1407 3218
rect 1473 1218 1503 3218
rect 1569 1218 1599 3218
rect 1665 1218 1695 3218
rect 1761 1218 1791 3218
rect 1857 1218 1887 3218
rect 1953 1218 1983 3218
rect 2049 1218 2079 3218
rect 2145 1218 2175 3218
rect 2241 1218 2271 3218
rect 2337 1218 2367 3218
rect 2433 1218 2463 3218
rect 2529 1218 2559 3218
rect 2625 1218 2655 3218
rect 2721 1218 2751 3218
rect 2817 1218 2847 3218
rect -2847 -1000 -2817 1000
rect -2751 -1000 -2721 1000
rect -2655 -1000 -2625 1000
rect -2559 -1000 -2529 1000
rect -2463 -1000 -2433 1000
rect -2367 -1000 -2337 1000
rect -2271 -1000 -2241 1000
rect -2175 -1000 -2145 1000
rect -2079 -1000 -2049 1000
rect -1983 -1000 -1953 1000
rect -1887 -1000 -1857 1000
rect -1791 -1000 -1761 1000
rect -1695 -1000 -1665 1000
rect -1599 -1000 -1569 1000
rect -1503 -1000 -1473 1000
rect -1407 -1000 -1377 1000
rect -1311 -1000 -1281 1000
rect -1215 -1000 -1185 1000
rect -1119 -1000 -1089 1000
rect -1023 -1000 -993 1000
rect -927 -1000 -897 1000
rect -831 -1000 -801 1000
rect -735 -1000 -705 1000
rect -639 -1000 -609 1000
rect -543 -1000 -513 1000
rect -447 -1000 -417 1000
rect -351 -1000 -321 1000
rect -255 -1000 -225 1000
rect -159 -1000 -129 1000
rect -63 -1000 -33 1000
rect 33 -1000 63 1000
rect 129 -1000 159 1000
rect 225 -1000 255 1000
rect 321 -1000 351 1000
rect 417 -1000 447 1000
rect 513 -1000 543 1000
rect 609 -1000 639 1000
rect 705 -1000 735 1000
rect 801 -1000 831 1000
rect 897 -1000 927 1000
rect 993 -1000 1023 1000
rect 1089 -1000 1119 1000
rect 1185 -1000 1215 1000
rect 1281 -1000 1311 1000
rect 1377 -1000 1407 1000
rect 1473 -1000 1503 1000
rect 1569 -1000 1599 1000
rect 1665 -1000 1695 1000
rect 1761 -1000 1791 1000
rect 1857 -1000 1887 1000
rect 1953 -1000 1983 1000
rect 2049 -1000 2079 1000
rect 2145 -1000 2175 1000
rect 2241 -1000 2271 1000
rect 2337 -1000 2367 1000
rect 2433 -1000 2463 1000
rect 2529 -1000 2559 1000
rect 2625 -1000 2655 1000
rect 2721 -1000 2751 1000
rect 2817 -1000 2847 1000
rect -2847 -3218 -2817 -1218
rect -2751 -3218 -2721 -1218
rect -2655 -3218 -2625 -1218
rect -2559 -3218 -2529 -1218
rect -2463 -3218 -2433 -1218
rect -2367 -3218 -2337 -1218
rect -2271 -3218 -2241 -1218
rect -2175 -3218 -2145 -1218
rect -2079 -3218 -2049 -1218
rect -1983 -3218 -1953 -1218
rect -1887 -3218 -1857 -1218
rect -1791 -3218 -1761 -1218
rect -1695 -3218 -1665 -1218
rect -1599 -3218 -1569 -1218
rect -1503 -3218 -1473 -1218
rect -1407 -3218 -1377 -1218
rect -1311 -3218 -1281 -1218
rect -1215 -3218 -1185 -1218
rect -1119 -3218 -1089 -1218
rect -1023 -3218 -993 -1218
rect -927 -3218 -897 -1218
rect -831 -3218 -801 -1218
rect -735 -3218 -705 -1218
rect -639 -3218 -609 -1218
rect -543 -3218 -513 -1218
rect -447 -3218 -417 -1218
rect -351 -3218 -321 -1218
rect -255 -3218 -225 -1218
rect -159 -3218 -129 -1218
rect -63 -3218 -33 -1218
rect 33 -3218 63 -1218
rect 129 -3218 159 -1218
rect 225 -3218 255 -1218
rect 321 -3218 351 -1218
rect 417 -3218 447 -1218
rect 513 -3218 543 -1218
rect 609 -3218 639 -1218
rect 705 -3218 735 -1218
rect 801 -3218 831 -1218
rect 897 -3218 927 -1218
rect 993 -3218 1023 -1218
rect 1089 -3218 1119 -1218
rect 1185 -3218 1215 -1218
rect 1281 -3218 1311 -1218
rect 1377 -3218 1407 -1218
rect 1473 -3218 1503 -1218
rect 1569 -3218 1599 -1218
rect 1665 -3218 1695 -1218
rect 1761 -3218 1791 -1218
rect 1857 -3218 1887 -1218
rect 1953 -3218 1983 -1218
rect 2049 -3218 2079 -1218
rect 2145 -3218 2175 -1218
rect 2241 -3218 2271 -1218
rect 2337 -3218 2367 -1218
rect 2433 -3218 2463 -1218
rect 2529 -3218 2559 -1218
rect 2625 -3218 2655 -1218
rect 2721 -3218 2751 -1218
rect 2817 -3218 2847 -1218
<< ndiff >>
rect -2909 3206 -2847 3218
rect -2909 1230 -2897 3206
rect -2863 1230 -2847 3206
rect -2909 1218 -2847 1230
rect -2817 3206 -2751 3218
rect -2817 1230 -2801 3206
rect -2767 1230 -2751 3206
rect -2817 1218 -2751 1230
rect -2721 3206 -2655 3218
rect -2721 1230 -2705 3206
rect -2671 1230 -2655 3206
rect -2721 1218 -2655 1230
rect -2625 3206 -2559 3218
rect -2625 1230 -2609 3206
rect -2575 1230 -2559 3206
rect -2625 1218 -2559 1230
rect -2529 3206 -2463 3218
rect -2529 1230 -2513 3206
rect -2479 1230 -2463 3206
rect -2529 1218 -2463 1230
rect -2433 3206 -2367 3218
rect -2433 1230 -2417 3206
rect -2383 1230 -2367 3206
rect -2433 1218 -2367 1230
rect -2337 3206 -2271 3218
rect -2337 1230 -2321 3206
rect -2287 1230 -2271 3206
rect -2337 1218 -2271 1230
rect -2241 3206 -2175 3218
rect -2241 1230 -2225 3206
rect -2191 1230 -2175 3206
rect -2241 1218 -2175 1230
rect -2145 3206 -2079 3218
rect -2145 1230 -2129 3206
rect -2095 1230 -2079 3206
rect -2145 1218 -2079 1230
rect -2049 3206 -1983 3218
rect -2049 1230 -2033 3206
rect -1999 1230 -1983 3206
rect -2049 1218 -1983 1230
rect -1953 3206 -1887 3218
rect -1953 1230 -1937 3206
rect -1903 1230 -1887 3206
rect -1953 1218 -1887 1230
rect -1857 3206 -1791 3218
rect -1857 1230 -1841 3206
rect -1807 1230 -1791 3206
rect -1857 1218 -1791 1230
rect -1761 3206 -1695 3218
rect -1761 1230 -1745 3206
rect -1711 1230 -1695 3206
rect -1761 1218 -1695 1230
rect -1665 3206 -1599 3218
rect -1665 1230 -1649 3206
rect -1615 1230 -1599 3206
rect -1665 1218 -1599 1230
rect -1569 3206 -1503 3218
rect -1569 1230 -1553 3206
rect -1519 1230 -1503 3206
rect -1569 1218 -1503 1230
rect -1473 3206 -1407 3218
rect -1473 1230 -1457 3206
rect -1423 1230 -1407 3206
rect -1473 1218 -1407 1230
rect -1377 3206 -1311 3218
rect -1377 1230 -1361 3206
rect -1327 1230 -1311 3206
rect -1377 1218 -1311 1230
rect -1281 3206 -1215 3218
rect -1281 1230 -1265 3206
rect -1231 1230 -1215 3206
rect -1281 1218 -1215 1230
rect -1185 3206 -1119 3218
rect -1185 1230 -1169 3206
rect -1135 1230 -1119 3206
rect -1185 1218 -1119 1230
rect -1089 3206 -1023 3218
rect -1089 1230 -1073 3206
rect -1039 1230 -1023 3206
rect -1089 1218 -1023 1230
rect -993 3206 -927 3218
rect -993 1230 -977 3206
rect -943 1230 -927 3206
rect -993 1218 -927 1230
rect -897 3206 -831 3218
rect -897 1230 -881 3206
rect -847 1230 -831 3206
rect -897 1218 -831 1230
rect -801 3206 -735 3218
rect -801 1230 -785 3206
rect -751 1230 -735 3206
rect -801 1218 -735 1230
rect -705 3206 -639 3218
rect -705 1230 -689 3206
rect -655 1230 -639 3206
rect -705 1218 -639 1230
rect -609 3206 -543 3218
rect -609 1230 -593 3206
rect -559 1230 -543 3206
rect -609 1218 -543 1230
rect -513 3206 -447 3218
rect -513 1230 -497 3206
rect -463 1230 -447 3206
rect -513 1218 -447 1230
rect -417 3206 -351 3218
rect -417 1230 -401 3206
rect -367 1230 -351 3206
rect -417 1218 -351 1230
rect -321 3206 -255 3218
rect -321 1230 -305 3206
rect -271 1230 -255 3206
rect -321 1218 -255 1230
rect -225 3206 -159 3218
rect -225 1230 -209 3206
rect -175 1230 -159 3206
rect -225 1218 -159 1230
rect -129 3206 -63 3218
rect -129 1230 -113 3206
rect -79 1230 -63 3206
rect -129 1218 -63 1230
rect -33 3206 33 3218
rect -33 1230 -17 3206
rect 17 1230 33 3206
rect -33 1218 33 1230
rect 63 3206 129 3218
rect 63 1230 79 3206
rect 113 1230 129 3206
rect 63 1218 129 1230
rect 159 3206 225 3218
rect 159 1230 175 3206
rect 209 1230 225 3206
rect 159 1218 225 1230
rect 255 3206 321 3218
rect 255 1230 271 3206
rect 305 1230 321 3206
rect 255 1218 321 1230
rect 351 3206 417 3218
rect 351 1230 367 3206
rect 401 1230 417 3206
rect 351 1218 417 1230
rect 447 3206 513 3218
rect 447 1230 463 3206
rect 497 1230 513 3206
rect 447 1218 513 1230
rect 543 3206 609 3218
rect 543 1230 559 3206
rect 593 1230 609 3206
rect 543 1218 609 1230
rect 639 3206 705 3218
rect 639 1230 655 3206
rect 689 1230 705 3206
rect 639 1218 705 1230
rect 735 3206 801 3218
rect 735 1230 751 3206
rect 785 1230 801 3206
rect 735 1218 801 1230
rect 831 3206 897 3218
rect 831 1230 847 3206
rect 881 1230 897 3206
rect 831 1218 897 1230
rect 927 3206 993 3218
rect 927 1230 943 3206
rect 977 1230 993 3206
rect 927 1218 993 1230
rect 1023 3206 1089 3218
rect 1023 1230 1039 3206
rect 1073 1230 1089 3206
rect 1023 1218 1089 1230
rect 1119 3206 1185 3218
rect 1119 1230 1135 3206
rect 1169 1230 1185 3206
rect 1119 1218 1185 1230
rect 1215 3206 1281 3218
rect 1215 1230 1231 3206
rect 1265 1230 1281 3206
rect 1215 1218 1281 1230
rect 1311 3206 1377 3218
rect 1311 1230 1327 3206
rect 1361 1230 1377 3206
rect 1311 1218 1377 1230
rect 1407 3206 1473 3218
rect 1407 1230 1423 3206
rect 1457 1230 1473 3206
rect 1407 1218 1473 1230
rect 1503 3206 1569 3218
rect 1503 1230 1519 3206
rect 1553 1230 1569 3206
rect 1503 1218 1569 1230
rect 1599 3206 1665 3218
rect 1599 1230 1615 3206
rect 1649 1230 1665 3206
rect 1599 1218 1665 1230
rect 1695 3206 1761 3218
rect 1695 1230 1711 3206
rect 1745 1230 1761 3206
rect 1695 1218 1761 1230
rect 1791 3206 1857 3218
rect 1791 1230 1807 3206
rect 1841 1230 1857 3206
rect 1791 1218 1857 1230
rect 1887 3206 1953 3218
rect 1887 1230 1903 3206
rect 1937 1230 1953 3206
rect 1887 1218 1953 1230
rect 1983 3206 2049 3218
rect 1983 1230 1999 3206
rect 2033 1230 2049 3206
rect 1983 1218 2049 1230
rect 2079 3206 2145 3218
rect 2079 1230 2095 3206
rect 2129 1230 2145 3206
rect 2079 1218 2145 1230
rect 2175 3206 2241 3218
rect 2175 1230 2191 3206
rect 2225 1230 2241 3206
rect 2175 1218 2241 1230
rect 2271 3206 2337 3218
rect 2271 1230 2287 3206
rect 2321 1230 2337 3206
rect 2271 1218 2337 1230
rect 2367 3206 2433 3218
rect 2367 1230 2383 3206
rect 2417 1230 2433 3206
rect 2367 1218 2433 1230
rect 2463 3206 2529 3218
rect 2463 1230 2479 3206
rect 2513 1230 2529 3206
rect 2463 1218 2529 1230
rect 2559 3206 2625 3218
rect 2559 1230 2575 3206
rect 2609 1230 2625 3206
rect 2559 1218 2625 1230
rect 2655 3206 2721 3218
rect 2655 1230 2671 3206
rect 2705 1230 2721 3206
rect 2655 1218 2721 1230
rect 2751 3206 2817 3218
rect 2751 1230 2767 3206
rect 2801 1230 2817 3206
rect 2751 1218 2817 1230
rect 2847 3206 2909 3218
rect 2847 1230 2863 3206
rect 2897 1230 2909 3206
rect 2847 1218 2909 1230
rect -2909 988 -2847 1000
rect -2909 -988 -2897 988
rect -2863 -988 -2847 988
rect -2909 -1000 -2847 -988
rect -2817 988 -2751 1000
rect -2817 -988 -2801 988
rect -2767 -988 -2751 988
rect -2817 -1000 -2751 -988
rect -2721 988 -2655 1000
rect -2721 -988 -2705 988
rect -2671 -988 -2655 988
rect -2721 -1000 -2655 -988
rect -2625 988 -2559 1000
rect -2625 -988 -2609 988
rect -2575 -988 -2559 988
rect -2625 -1000 -2559 -988
rect -2529 988 -2463 1000
rect -2529 -988 -2513 988
rect -2479 -988 -2463 988
rect -2529 -1000 -2463 -988
rect -2433 988 -2367 1000
rect -2433 -988 -2417 988
rect -2383 -988 -2367 988
rect -2433 -1000 -2367 -988
rect -2337 988 -2271 1000
rect -2337 -988 -2321 988
rect -2287 -988 -2271 988
rect -2337 -1000 -2271 -988
rect -2241 988 -2175 1000
rect -2241 -988 -2225 988
rect -2191 -988 -2175 988
rect -2241 -1000 -2175 -988
rect -2145 988 -2079 1000
rect -2145 -988 -2129 988
rect -2095 -988 -2079 988
rect -2145 -1000 -2079 -988
rect -2049 988 -1983 1000
rect -2049 -988 -2033 988
rect -1999 -988 -1983 988
rect -2049 -1000 -1983 -988
rect -1953 988 -1887 1000
rect -1953 -988 -1937 988
rect -1903 -988 -1887 988
rect -1953 -1000 -1887 -988
rect -1857 988 -1791 1000
rect -1857 -988 -1841 988
rect -1807 -988 -1791 988
rect -1857 -1000 -1791 -988
rect -1761 988 -1695 1000
rect -1761 -988 -1745 988
rect -1711 -988 -1695 988
rect -1761 -1000 -1695 -988
rect -1665 988 -1599 1000
rect -1665 -988 -1649 988
rect -1615 -988 -1599 988
rect -1665 -1000 -1599 -988
rect -1569 988 -1503 1000
rect -1569 -988 -1553 988
rect -1519 -988 -1503 988
rect -1569 -1000 -1503 -988
rect -1473 988 -1407 1000
rect -1473 -988 -1457 988
rect -1423 -988 -1407 988
rect -1473 -1000 -1407 -988
rect -1377 988 -1311 1000
rect -1377 -988 -1361 988
rect -1327 -988 -1311 988
rect -1377 -1000 -1311 -988
rect -1281 988 -1215 1000
rect -1281 -988 -1265 988
rect -1231 -988 -1215 988
rect -1281 -1000 -1215 -988
rect -1185 988 -1119 1000
rect -1185 -988 -1169 988
rect -1135 -988 -1119 988
rect -1185 -1000 -1119 -988
rect -1089 988 -1023 1000
rect -1089 -988 -1073 988
rect -1039 -988 -1023 988
rect -1089 -1000 -1023 -988
rect -993 988 -927 1000
rect -993 -988 -977 988
rect -943 -988 -927 988
rect -993 -1000 -927 -988
rect -897 988 -831 1000
rect -897 -988 -881 988
rect -847 -988 -831 988
rect -897 -1000 -831 -988
rect -801 988 -735 1000
rect -801 -988 -785 988
rect -751 -988 -735 988
rect -801 -1000 -735 -988
rect -705 988 -639 1000
rect -705 -988 -689 988
rect -655 -988 -639 988
rect -705 -1000 -639 -988
rect -609 988 -543 1000
rect -609 -988 -593 988
rect -559 -988 -543 988
rect -609 -1000 -543 -988
rect -513 988 -447 1000
rect -513 -988 -497 988
rect -463 -988 -447 988
rect -513 -1000 -447 -988
rect -417 988 -351 1000
rect -417 -988 -401 988
rect -367 -988 -351 988
rect -417 -1000 -351 -988
rect -321 988 -255 1000
rect -321 -988 -305 988
rect -271 -988 -255 988
rect -321 -1000 -255 -988
rect -225 988 -159 1000
rect -225 -988 -209 988
rect -175 -988 -159 988
rect -225 -1000 -159 -988
rect -129 988 -63 1000
rect -129 -988 -113 988
rect -79 -988 -63 988
rect -129 -1000 -63 -988
rect -33 988 33 1000
rect -33 -988 -17 988
rect 17 -988 33 988
rect -33 -1000 33 -988
rect 63 988 129 1000
rect 63 -988 79 988
rect 113 -988 129 988
rect 63 -1000 129 -988
rect 159 988 225 1000
rect 159 -988 175 988
rect 209 -988 225 988
rect 159 -1000 225 -988
rect 255 988 321 1000
rect 255 -988 271 988
rect 305 -988 321 988
rect 255 -1000 321 -988
rect 351 988 417 1000
rect 351 -988 367 988
rect 401 -988 417 988
rect 351 -1000 417 -988
rect 447 988 513 1000
rect 447 -988 463 988
rect 497 -988 513 988
rect 447 -1000 513 -988
rect 543 988 609 1000
rect 543 -988 559 988
rect 593 -988 609 988
rect 543 -1000 609 -988
rect 639 988 705 1000
rect 639 -988 655 988
rect 689 -988 705 988
rect 639 -1000 705 -988
rect 735 988 801 1000
rect 735 -988 751 988
rect 785 -988 801 988
rect 735 -1000 801 -988
rect 831 988 897 1000
rect 831 -988 847 988
rect 881 -988 897 988
rect 831 -1000 897 -988
rect 927 988 993 1000
rect 927 -988 943 988
rect 977 -988 993 988
rect 927 -1000 993 -988
rect 1023 988 1089 1000
rect 1023 -988 1039 988
rect 1073 -988 1089 988
rect 1023 -1000 1089 -988
rect 1119 988 1185 1000
rect 1119 -988 1135 988
rect 1169 -988 1185 988
rect 1119 -1000 1185 -988
rect 1215 988 1281 1000
rect 1215 -988 1231 988
rect 1265 -988 1281 988
rect 1215 -1000 1281 -988
rect 1311 988 1377 1000
rect 1311 -988 1327 988
rect 1361 -988 1377 988
rect 1311 -1000 1377 -988
rect 1407 988 1473 1000
rect 1407 -988 1423 988
rect 1457 -988 1473 988
rect 1407 -1000 1473 -988
rect 1503 988 1569 1000
rect 1503 -988 1519 988
rect 1553 -988 1569 988
rect 1503 -1000 1569 -988
rect 1599 988 1665 1000
rect 1599 -988 1615 988
rect 1649 -988 1665 988
rect 1599 -1000 1665 -988
rect 1695 988 1761 1000
rect 1695 -988 1711 988
rect 1745 -988 1761 988
rect 1695 -1000 1761 -988
rect 1791 988 1857 1000
rect 1791 -988 1807 988
rect 1841 -988 1857 988
rect 1791 -1000 1857 -988
rect 1887 988 1953 1000
rect 1887 -988 1903 988
rect 1937 -988 1953 988
rect 1887 -1000 1953 -988
rect 1983 988 2049 1000
rect 1983 -988 1999 988
rect 2033 -988 2049 988
rect 1983 -1000 2049 -988
rect 2079 988 2145 1000
rect 2079 -988 2095 988
rect 2129 -988 2145 988
rect 2079 -1000 2145 -988
rect 2175 988 2241 1000
rect 2175 -988 2191 988
rect 2225 -988 2241 988
rect 2175 -1000 2241 -988
rect 2271 988 2337 1000
rect 2271 -988 2287 988
rect 2321 -988 2337 988
rect 2271 -1000 2337 -988
rect 2367 988 2433 1000
rect 2367 -988 2383 988
rect 2417 -988 2433 988
rect 2367 -1000 2433 -988
rect 2463 988 2529 1000
rect 2463 -988 2479 988
rect 2513 -988 2529 988
rect 2463 -1000 2529 -988
rect 2559 988 2625 1000
rect 2559 -988 2575 988
rect 2609 -988 2625 988
rect 2559 -1000 2625 -988
rect 2655 988 2721 1000
rect 2655 -988 2671 988
rect 2705 -988 2721 988
rect 2655 -1000 2721 -988
rect 2751 988 2817 1000
rect 2751 -988 2767 988
rect 2801 -988 2817 988
rect 2751 -1000 2817 -988
rect 2847 988 2909 1000
rect 2847 -988 2863 988
rect 2897 -988 2909 988
rect 2847 -1000 2909 -988
rect -2909 -1230 -2847 -1218
rect -2909 -3206 -2897 -1230
rect -2863 -3206 -2847 -1230
rect -2909 -3218 -2847 -3206
rect -2817 -1230 -2751 -1218
rect -2817 -3206 -2801 -1230
rect -2767 -3206 -2751 -1230
rect -2817 -3218 -2751 -3206
rect -2721 -1230 -2655 -1218
rect -2721 -3206 -2705 -1230
rect -2671 -3206 -2655 -1230
rect -2721 -3218 -2655 -3206
rect -2625 -1230 -2559 -1218
rect -2625 -3206 -2609 -1230
rect -2575 -3206 -2559 -1230
rect -2625 -3218 -2559 -3206
rect -2529 -1230 -2463 -1218
rect -2529 -3206 -2513 -1230
rect -2479 -3206 -2463 -1230
rect -2529 -3218 -2463 -3206
rect -2433 -1230 -2367 -1218
rect -2433 -3206 -2417 -1230
rect -2383 -3206 -2367 -1230
rect -2433 -3218 -2367 -3206
rect -2337 -1230 -2271 -1218
rect -2337 -3206 -2321 -1230
rect -2287 -3206 -2271 -1230
rect -2337 -3218 -2271 -3206
rect -2241 -1230 -2175 -1218
rect -2241 -3206 -2225 -1230
rect -2191 -3206 -2175 -1230
rect -2241 -3218 -2175 -3206
rect -2145 -1230 -2079 -1218
rect -2145 -3206 -2129 -1230
rect -2095 -3206 -2079 -1230
rect -2145 -3218 -2079 -3206
rect -2049 -1230 -1983 -1218
rect -2049 -3206 -2033 -1230
rect -1999 -3206 -1983 -1230
rect -2049 -3218 -1983 -3206
rect -1953 -1230 -1887 -1218
rect -1953 -3206 -1937 -1230
rect -1903 -3206 -1887 -1230
rect -1953 -3218 -1887 -3206
rect -1857 -1230 -1791 -1218
rect -1857 -3206 -1841 -1230
rect -1807 -3206 -1791 -1230
rect -1857 -3218 -1791 -3206
rect -1761 -1230 -1695 -1218
rect -1761 -3206 -1745 -1230
rect -1711 -3206 -1695 -1230
rect -1761 -3218 -1695 -3206
rect -1665 -1230 -1599 -1218
rect -1665 -3206 -1649 -1230
rect -1615 -3206 -1599 -1230
rect -1665 -3218 -1599 -3206
rect -1569 -1230 -1503 -1218
rect -1569 -3206 -1553 -1230
rect -1519 -3206 -1503 -1230
rect -1569 -3218 -1503 -3206
rect -1473 -1230 -1407 -1218
rect -1473 -3206 -1457 -1230
rect -1423 -3206 -1407 -1230
rect -1473 -3218 -1407 -3206
rect -1377 -1230 -1311 -1218
rect -1377 -3206 -1361 -1230
rect -1327 -3206 -1311 -1230
rect -1377 -3218 -1311 -3206
rect -1281 -1230 -1215 -1218
rect -1281 -3206 -1265 -1230
rect -1231 -3206 -1215 -1230
rect -1281 -3218 -1215 -3206
rect -1185 -1230 -1119 -1218
rect -1185 -3206 -1169 -1230
rect -1135 -3206 -1119 -1230
rect -1185 -3218 -1119 -3206
rect -1089 -1230 -1023 -1218
rect -1089 -3206 -1073 -1230
rect -1039 -3206 -1023 -1230
rect -1089 -3218 -1023 -3206
rect -993 -1230 -927 -1218
rect -993 -3206 -977 -1230
rect -943 -3206 -927 -1230
rect -993 -3218 -927 -3206
rect -897 -1230 -831 -1218
rect -897 -3206 -881 -1230
rect -847 -3206 -831 -1230
rect -897 -3218 -831 -3206
rect -801 -1230 -735 -1218
rect -801 -3206 -785 -1230
rect -751 -3206 -735 -1230
rect -801 -3218 -735 -3206
rect -705 -1230 -639 -1218
rect -705 -3206 -689 -1230
rect -655 -3206 -639 -1230
rect -705 -3218 -639 -3206
rect -609 -1230 -543 -1218
rect -609 -3206 -593 -1230
rect -559 -3206 -543 -1230
rect -609 -3218 -543 -3206
rect -513 -1230 -447 -1218
rect -513 -3206 -497 -1230
rect -463 -3206 -447 -1230
rect -513 -3218 -447 -3206
rect -417 -1230 -351 -1218
rect -417 -3206 -401 -1230
rect -367 -3206 -351 -1230
rect -417 -3218 -351 -3206
rect -321 -1230 -255 -1218
rect -321 -3206 -305 -1230
rect -271 -3206 -255 -1230
rect -321 -3218 -255 -3206
rect -225 -1230 -159 -1218
rect -225 -3206 -209 -1230
rect -175 -3206 -159 -1230
rect -225 -3218 -159 -3206
rect -129 -1230 -63 -1218
rect -129 -3206 -113 -1230
rect -79 -3206 -63 -1230
rect -129 -3218 -63 -3206
rect -33 -1230 33 -1218
rect -33 -3206 -17 -1230
rect 17 -3206 33 -1230
rect -33 -3218 33 -3206
rect 63 -1230 129 -1218
rect 63 -3206 79 -1230
rect 113 -3206 129 -1230
rect 63 -3218 129 -3206
rect 159 -1230 225 -1218
rect 159 -3206 175 -1230
rect 209 -3206 225 -1230
rect 159 -3218 225 -3206
rect 255 -1230 321 -1218
rect 255 -3206 271 -1230
rect 305 -3206 321 -1230
rect 255 -3218 321 -3206
rect 351 -1230 417 -1218
rect 351 -3206 367 -1230
rect 401 -3206 417 -1230
rect 351 -3218 417 -3206
rect 447 -1230 513 -1218
rect 447 -3206 463 -1230
rect 497 -3206 513 -1230
rect 447 -3218 513 -3206
rect 543 -1230 609 -1218
rect 543 -3206 559 -1230
rect 593 -3206 609 -1230
rect 543 -3218 609 -3206
rect 639 -1230 705 -1218
rect 639 -3206 655 -1230
rect 689 -3206 705 -1230
rect 639 -3218 705 -3206
rect 735 -1230 801 -1218
rect 735 -3206 751 -1230
rect 785 -3206 801 -1230
rect 735 -3218 801 -3206
rect 831 -1230 897 -1218
rect 831 -3206 847 -1230
rect 881 -3206 897 -1230
rect 831 -3218 897 -3206
rect 927 -1230 993 -1218
rect 927 -3206 943 -1230
rect 977 -3206 993 -1230
rect 927 -3218 993 -3206
rect 1023 -1230 1089 -1218
rect 1023 -3206 1039 -1230
rect 1073 -3206 1089 -1230
rect 1023 -3218 1089 -3206
rect 1119 -1230 1185 -1218
rect 1119 -3206 1135 -1230
rect 1169 -3206 1185 -1230
rect 1119 -3218 1185 -3206
rect 1215 -1230 1281 -1218
rect 1215 -3206 1231 -1230
rect 1265 -3206 1281 -1230
rect 1215 -3218 1281 -3206
rect 1311 -1230 1377 -1218
rect 1311 -3206 1327 -1230
rect 1361 -3206 1377 -1230
rect 1311 -3218 1377 -3206
rect 1407 -1230 1473 -1218
rect 1407 -3206 1423 -1230
rect 1457 -3206 1473 -1230
rect 1407 -3218 1473 -3206
rect 1503 -1230 1569 -1218
rect 1503 -3206 1519 -1230
rect 1553 -3206 1569 -1230
rect 1503 -3218 1569 -3206
rect 1599 -1230 1665 -1218
rect 1599 -3206 1615 -1230
rect 1649 -3206 1665 -1230
rect 1599 -3218 1665 -3206
rect 1695 -1230 1761 -1218
rect 1695 -3206 1711 -1230
rect 1745 -3206 1761 -1230
rect 1695 -3218 1761 -3206
rect 1791 -1230 1857 -1218
rect 1791 -3206 1807 -1230
rect 1841 -3206 1857 -1230
rect 1791 -3218 1857 -3206
rect 1887 -1230 1953 -1218
rect 1887 -3206 1903 -1230
rect 1937 -3206 1953 -1230
rect 1887 -3218 1953 -3206
rect 1983 -1230 2049 -1218
rect 1983 -3206 1999 -1230
rect 2033 -3206 2049 -1230
rect 1983 -3218 2049 -3206
rect 2079 -1230 2145 -1218
rect 2079 -3206 2095 -1230
rect 2129 -3206 2145 -1230
rect 2079 -3218 2145 -3206
rect 2175 -1230 2241 -1218
rect 2175 -3206 2191 -1230
rect 2225 -3206 2241 -1230
rect 2175 -3218 2241 -3206
rect 2271 -1230 2337 -1218
rect 2271 -3206 2287 -1230
rect 2321 -3206 2337 -1230
rect 2271 -3218 2337 -3206
rect 2367 -1230 2433 -1218
rect 2367 -3206 2383 -1230
rect 2417 -3206 2433 -1230
rect 2367 -3218 2433 -3206
rect 2463 -1230 2529 -1218
rect 2463 -3206 2479 -1230
rect 2513 -3206 2529 -1230
rect 2463 -3218 2529 -3206
rect 2559 -1230 2625 -1218
rect 2559 -3206 2575 -1230
rect 2609 -3206 2625 -1230
rect 2559 -3218 2625 -3206
rect 2655 -1230 2721 -1218
rect 2655 -3206 2671 -1230
rect 2705 -3206 2721 -1230
rect 2655 -3218 2721 -3206
rect 2751 -1230 2817 -1218
rect 2751 -3206 2767 -1230
rect 2801 -3206 2817 -1230
rect 2751 -3218 2817 -3206
rect 2847 -1230 2909 -1218
rect 2847 -3206 2863 -1230
rect 2897 -3206 2909 -1230
rect 2847 -3218 2909 -3206
<< ndiffc >>
rect -2897 1230 -2863 3206
rect -2801 1230 -2767 3206
rect -2705 1230 -2671 3206
rect -2609 1230 -2575 3206
rect -2513 1230 -2479 3206
rect -2417 1230 -2383 3206
rect -2321 1230 -2287 3206
rect -2225 1230 -2191 3206
rect -2129 1230 -2095 3206
rect -2033 1230 -1999 3206
rect -1937 1230 -1903 3206
rect -1841 1230 -1807 3206
rect -1745 1230 -1711 3206
rect -1649 1230 -1615 3206
rect -1553 1230 -1519 3206
rect -1457 1230 -1423 3206
rect -1361 1230 -1327 3206
rect -1265 1230 -1231 3206
rect -1169 1230 -1135 3206
rect -1073 1230 -1039 3206
rect -977 1230 -943 3206
rect -881 1230 -847 3206
rect -785 1230 -751 3206
rect -689 1230 -655 3206
rect -593 1230 -559 3206
rect -497 1230 -463 3206
rect -401 1230 -367 3206
rect -305 1230 -271 3206
rect -209 1230 -175 3206
rect -113 1230 -79 3206
rect -17 1230 17 3206
rect 79 1230 113 3206
rect 175 1230 209 3206
rect 271 1230 305 3206
rect 367 1230 401 3206
rect 463 1230 497 3206
rect 559 1230 593 3206
rect 655 1230 689 3206
rect 751 1230 785 3206
rect 847 1230 881 3206
rect 943 1230 977 3206
rect 1039 1230 1073 3206
rect 1135 1230 1169 3206
rect 1231 1230 1265 3206
rect 1327 1230 1361 3206
rect 1423 1230 1457 3206
rect 1519 1230 1553 3206
rect 1615 1230 1649 3206
rect 1711 1230 1745 3206
rect 1807 1230 1841 3206
rect 1903 1230 1937 3206
rect 1999 1230 2033 3206
rect 2095 1230 2129 3206
rect 2191 1230 2225 3206
rect 2287 1230 2321 3206
rect 2383 1230 2417 3206
rect 2479 1230 2513 3206
rect 2575 1230 2609 3206
rect 2671 1230 2705 3206
rect 2767 1230 2801 3206
rect 2863 1230 2897 3206
rect -2897 -988 -2863 988
rect -2801 -988 -2767 988
rect -2705 -988 -2671 988
rect -2609 -988 -2575 988
rect -2513 -988 -2479 988
rect -2417 -988 -2383 988
rect -2321 -988 -2287 988
rect -2225 -988 -2191 988
rect -2129 -988 -2095 988
rect -2033 -988 -1999 988
rect -1937 -988 -1903 988
rect -1841 -988 -1807 988
rect -1745 -988 -1711 988
rect -1649 -988 -1615 988
rect -1553 -988 -1519 988
rect -1457 -988 -1423 988
rect -1361 -988 -1327 988
rect -1265 -988 -1231 988
rect -1169 -988 -1135 988
rect -1073 -988 -1039 988
rect -977 -988 -943 988
rect -881 -988 -847 988
rect -785 -988 -751 988
rect -689 -988 -655 988
rect -593 -988 -559 988
rect -497 -988 -463 988
rect -401 -988 -367 988
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect 367 -988 401 988
rect 463 -988 497 988
rect 559 -988 593 988
rect 655 -988 689 988
rect 751 -988 785 988
rect 847 -988 881 988
rect 943 -988 977 988
rect 1039 -988 1073 988
rect 1135 -988 1169 988
rect 1231 -988 1265 988
rect 1327 -988 1361 988
rect 1423 -988 1457 988
rect 1519 -988 1553 988
rect 1615 -988 1649 988
rect 1711 -988 1745 988
rect 1807 -988 1841 988
rect 1903 -988 1937 988
rect 1999 -988 2033 988
rect 2095 -988 2129 988
rect 2191 -988 2225 988
rect 2287 -988 2321 988
rect 2383 -988 2417 988
rect 2479 -988 2513 988
rect 2575 -988 2609 988
rect 2671 -988 2705 988
rect 2767 -988 2801 988
rect 2863 -988 2897 988
rect -2897 -3206 -2863 -1230
rect -2801 -3206 -2767 -1230
rect -2705 -3206 -2671 -1230
rect -2609 -3206 -2575 -1230
rect -2513 -3206 -2479 -1230
rect -2417 -3206 -2383 -1230
rect -2321 -3206 -2287 -1230
rect -2225 -3206 -2191 -1230
rect -2129 -3206 -2095 -1230
rect -2033 -3206 -1999 -1230
rect -1937 -3206 -1903 -1230
rect -1841 -3206 -1807 -1230
rect -1745 -3206 -1711 -1230
rect -1649 -3206 -1615 -1230
rect -1553 -3206 -1519 -1230
rect -1457 -3206 -1423 -1230
rect -1361 -3206 -1327 -1230
rect -1265 -3206 -1231 -1230
rect -1169 -3206 -1135 -1230
rect -1073 -3206 -1039 -1230
rect -977 -3206 -943 -1230
rect -881 -3206 -847 -1230
rect -785 -3206 -751 -1230
rect -689 -3206 -655 -1230
rect -593 -3206 -559 -1230
rect -497 -3206 -463 -1230
rect -401 -3206 -367 -1230
rect -305 -3206 -271 -1230
rect -209 -3206 -175 -1230
rect -113 -3206 -79 -1230
rect -17 -3206 17 -1230
rect 79 -3206 113 -1230
rect 175 -3206 209 -1230
rect 271 -3206 305 -1230
rect 367 -3206 401 -1230
rect 463 -3206 497 -1230
rect 559 -3206 593 -1230
rect 655 -3206 689 -1230
rect 751 -3206 785 -1230
rect 847 -3206 881 -1230
rect 943 -3206 977 -1230
rect 1039 -3206 1073 -1230
rect 1135 -3206 1169 -1230
rect 1231 -3206 1265 -1230
rect 1327 -3206 1361 -1230
rect 1423 -3206 1457 -1230
rect 1519 -3206 1553 -1230
rect 1615 -3206 1649 -1230
rect 1711 -3206 1745 -1230
rect 1807 -3206 1841 -1230
rect 1903 -3206 1937 -1230
rect 1999 -3206 2033 -1230
rect 2095 -3206 2129 -1230
rect 2191 -3206 2225 -1230
rect 2287 -3206 2321 -1230
rect 2383 -3206 2417 -1230
rect 2479 -3206 2513 -1230
rect 2575 -3206 2609 -1230
rect 2671 -3206 2705 -1230
rect 2767 -3206 2801 -1230
rect 2863 -3206 2897 -1230
<< poly >>
rect -2769 3290 -2703 3306
rect -2769 3256 -2753 3290
rect -2719 3256 -2703 3290
rect -2847 3218 -2817 3244
rect -2769 3240 -2703 3256
rect -2577 3290 -2511 3306
rect -2577 3256 -2561 3290
rect -2527 3256 -2511 3290
rect -2751 3218 -2721 3240
rect -2655 3218 -2625 3244
rect -2577 3240 -2511 3256
rect -2385 3290 -2319 3306
rect -2385 3256 -2369 3290
rect -2335 3256 -2319 3290
rect -2559 3218 -2529 3240
rect -2463 3218 -2433 3244
rect -2385 3240 -2319 3256
rect -2193 3290 -2127 3306
rect -2193 3256 -2177 3290
rect -2143 3256 -2127 3290
rect -2367 3218 -2337 3240
rect -2271 3218 -2241 3244
rect -2193 3240 -2127 3256
rect -2001 3290 -1935 3306
rect -2001 3256 -1985 3290
rect -1951 3256 -1935 3290
rect -2175 3218 -2145 3240
rect -2079 3218 -2049 3244
rect -2001 3240 -1935 3256
rect -1809 3290 -1743 3306
rect -1809 3256 -1793 3290
rect -1759 3256 -1743 3290
rect -1983 3218 -1953 3240
rect -1887 3218 -1857 3244
rect -1809 3240 -1743 3256
rect -1617 3290 -1551 3306
rect -1617 3256 -1601 3290
rect -1567 3256 -1551 3290
rect -1791 3218 -1761 3240
rect -1695 3218 -1665 3244
rect -1617 3240 -1551 3256
rect -1425 3290 -1359 3306
rect -1425 3256 -1409 3290
rect -1375 3256 -1359 3290
rect -1599 3218 -1569 3240
rect -1503 3218 -1473 3244
rect -1425 3240 -1359 3256
rect -1233 3290 -1167 3306
rect -1233 3256 -1217 3290
rect -1183 3256 -1167 3290
rect -1407 3218 -1377 3240
rect -1311 3218 -1281 3244
rect -1233 3240 -1167 3256
rect -1041 3290 -975 3306
rect -1041 3256 -1025 3290
rect -991 3256 -975 3290
rect -1215 3218 -1185 3240
rect -1119 3218 -1089 3244
rect -1041 3240 -975 3256
rect -849 3290 -783 3306
rect -849 3256 -833 3290
rect -799 3256 -783 3290
rect -1023 3218 -993 3240
rect -927 3218 -897 3244
rect -849 3240 -783 3256
rect -657 3290 -591 3306
rect -657 3256 -641 3290
rect -607 3256 -591 3290
rect -831 3218 -801 3240
rect -735 3218 -705 3244
rect -657 3240 -591 3256
rect -465 3290 -399 3306
rect -465 3256 -449 3290
rect -415 3256 -399 3290
rect -639 3218 -609 3240
rect -543 3218 -513 3244
rect -465 3240 -399 3256
rect -273 3290 -207 3306
rect -273 3256 -257 3290
rect -223 3256 -207 3290
rect -447 3218 -417 3240
rect -351 3218 -321 3244
rect -273 3240 -207 3256
rect -81 3290 -15 3306
rect -81 3256 -65 3290
rect -31 3256 -15 3290
rect -255 3218 -225 3240
rect -159 3218 -129 3244
rect -81 3240 -15 3256
rect 111 3290 177 3306
rect 111 3256 127 3290
rect 161 3256 177 3290
rect -63 3218 -33 3240
rect 33 3218 63 3244
rect 111 3240 177 3256
rect 303 3290 369 3306
rect 303 3256 319 3290
rect 353 3256 369 3290
rect 129 3218 159 3240
rect 225 3218 255 3244
rect 303 3240 369 3256
rect 495 3290 561 3306
rect 495 3256 511 3290
rect 545 3256 561 3290
rect 321 3218 351 3240
rect 417 3218 447 3244
rect 495 3240 561 3256
rect 687 3290 753 3306
rect 687 3256 703 3290
rect 737 3256 753 3290
rect 513 3218 543 3240
rect 609 3218 639 3244
rect 687 3240 753 3256
rect 879 3290 945 3306
rect 879 3256 895 3290
rect 929 3256 945 3290
rect 705 3218 735 3240
rect 801 3218 831 3244
rect 879 3240 945 3256
rect 1071 3290 1137 3306
rect 1071 3256 1087 3290
rect 1121 3256 1137 3290
rect 897 3218 927 3240
rect 993 3218 1023 3244
rect 1071 3240 1137 3256
rect 1263 3290 1329 3306
rect 1263 3256 1279 3290
rect 1313 3256 1329 3290
rect 1089 3218 1119 3240
rect 1185 3218 1215 3244
rect 1263 3240 1329 3256
rect 1455 3290 1521 3306
rect 1455 3256 1471 3290
rect 1505 3256 1521 3290
rect 1281 3218 1311 3240
rect 1377 3218 1407 3244
rect 1455 3240 1521 3256
rect 1647 3290 1713 3306
rect 1647 3256 1663 3290
rect 1697 3256 1713 3290
rect 1473 3218 1503 3240
rect 1569 3218 1599 3244
rect 1647 3240 1713 3256
rect 1839 3290 1905 3306
rect 1839 3256 1855 3290
rect 1889 3256 1905 3290
rect 1665 3218 1695 3240
rect 1761 3218 1791 3244
rect 1839 3240 1905 3256
rect 2031 3290 2097 3306
rect 2031 3256 2047 3290
rect 2081 3256 2097 3290
rect 1857 3218 1887 3240
rect 1953 3218 1983 3244
rect 2031 3240 2097 3256
rect 2223 3290 2289 3306
rect 2223 3256 2239 3290
rect 2273 3256 2289 3290
rect 2049 3218 2079 3240
rect 2145 3218 2175 3244
rect 2223 3240 2289 3256
rect 2415 3290 2481 3306
rect 2415 3256 2431 3290
rect 2465 3256 2481 3290
rect 2241 3218 2271 3240
rect 2337 3218 2367 3244
rect 2415 3240 2481 3256
rect 2607 3290 2673 3306
rect 2607 3256 2623 3290
rect 2657 3256 2673 3290
rect 2433 3218 2463 3240
rect 2529 3218 2559 3244
rect 2607 3240 2673 3256
rect 2799 3290 2865 3306
rect 2799 3256 2815 3290
rect 2849 3256 2865 3290
rect 2625 3218 2655 3240
rect 2721 3218 2751 3244
rect 2799 3240 2865 3256
rect 2817 3218 2847 3240
rect -2847 1196 -2817 1218
rect -2865 1180 -2799 1196
rect -2751 1192 -2721 1218
rect -2655 1196 -2625 1218
rect -2865 1146 -2849 1180
rect -2815 1146 -2799 1180
rect -2865 1130 -2799 1146
rect -2673 1180 -2607 1196
rect -2559 1192 -2529 1218
rect -2463 1196 -2433 1218
rect -2673 1146 -2657 1180
rect -2623 1146 -2607 1180
rect -2673 1130 -2607 1146
rect -2481 1180 -2415 1196
rect -2367 1192 -2337 1218
rect -2271 1196 -2241 1218
rect -2481 1146 -2465 1180
rect -2431 1146 -2415 1180
rect -2481 1130 -2415 1146
rect -2289 1180 -2223 1196
rect -2175 1192 -2145 1218
rect -2079 1196 -2049 1218
rect -2289 1146 -2273 1180
rect -2239 1146 -2223 1180
rect -2289 1130 -2223 1146
rect -2097 1180 -2031 1196
rect -1983 1192 -1953 1218
rect -1887 1196 -1857 1218
rect -2097 1146 -2081 1180
rect -2047 1146 -2031 1180
rect -2097 1130 -2031 1146
rect -1905 1180 -1839 1196
rect -1791 1192 -1761 1218
rect -1695 1196 -1665 1218
rect -1905 1146 -1889 1180
rect -1855 1146 -1839 1180
rect -1905 1130 -1839 1146
rect -1713 1180 -1647 1196
rect -1599 1192 -1569 1218
rect -1503 1196 -1473 1218
rect -1713 1146 -1697 1180
rect -1663 1146 -1647 1180
rect -1713 1130 -1647 1146
rect -1521 1180 -1455 1196
rect -1407 1192 -1377 1218
rect -1311 1196 -1281 1218
rect -1521 1146 -1505 1180
rect -1471 1146 -1455 1180
rect -1521 1130 -1455 1146
rect -1329 1180 -1263 1196
rect -1215 1192 -1185 1218
rect -1119 1196 -1089 1218
rect -1329 1146 -1313 1180
rect -1279 1146 -1263 1180
rect -1329 1130 -1263 1146
rect -1137 1180 -1071 1196
rect -1023 1192 -993 1218
rect -927 1196 -897 1218
rect -1137 1146 -1121 1180
rect -1087 1146 -1071 1180
rect -1137 1130 -1071 1146
rect -945 1180 -879 1196
rect -831 1192 -801 1218
rect -735 1196 -705 1218
rect -945 1146 -929 1180
rect -895 1146 -879 1180
rect -945 1130 -879 1146
rect -753 1180 -687 1196
rect -639 1192 -609 1218
rect -543 1196 -513 1218
rect -753 1146 -737 1180
rect -703 1146 -687 1180
rect -753 1130 -687 1146
rect -561 1180 -495 1196
rect -447 1192 -417 1218
rect -351 1196 -321 1218
rect -561 1146 -545 1180
rect -511 1146 -495 1180
rect -561 1130 -495 1146
rect -369 1180 -303 1196
rect -255 1192 -225 1218
rect -159 1196 -129 1218
rect -369 1146 -353 1180
rect -319 1146 -303 1180
rect -369 1130 -303 1146
rect -177 1180 -111 1196
rect -63 1192 -33 1218
rect 33 1196 63 1218
rect -177 1146 -161 1180
rect -127 1146 -111 1180
rect -177 1130 -111 1146
rect 15 1180 81 1196
rect 129 1192 159 1218
rect 225 1196 255 1218
rect 15 1146 31 1180
rect 65 1146 81 1180
rect 15 1130 81 1146
rect 207 1180 273 1196
rect 321 1192 351 1218
rect 417 1196 447 1218
rect 207 1146 223 1180
rect 257 1146 273 1180
rect 207 1130 273 1146
rect 399 1180 465 1196
rect 513 1192 543 1218
rect 609 1196 639 1218
rect 399 1146 415 1180
rect 449 1146 465 1180
rect 399 1130 465 1146
rect 591 1180 657 1196
rect 705 1192 735 1218
rect 801 1196 831 1218
rect 591 1146 607 1180
rect 641 1146 657 1180
rect 591 1130 657 1146
rect 783 1180 849 1196
rect 897 1192 927 1218
rect 993 1196 1023 1218
rect 783 1146 799 1180
rect 833 1146 849 1180
rect 783 1130 849 1146
rect 975 1180 1041 1196
rect 1089 1192 1119 1218
rect 1185 1196 1215 1218
rect 975 1146 991 1180
rect 1025 1146 1041 1180
rect 975 1130 1041 1146
rect 1167 1180 1233 1196
rect 1281 1192 1311 1218
rect 1377 1196 1407 1218
rect 1167 1146 1183 1180
rect 1217 1146 1233 1180
rect 1167 1130 1233 1146
rect 1359 1180 1425 1196
rect 1473 1192 1503 1218
rect 1569 1196 1599 1218
rect 1359 1146 1375 1180
rect 1409 1146 1425 1180
rect 1359 1130 1425 1146
rect 1551 1180 1617 1196
rect 1665 1192 1695 1218
rect 1761 1196 1791 1218
rect 1551 1146 1567 1180
rect 1601 1146 1617 1180
rect 1551 1130 1617 1146
rect 1743 1180 1809 1196
rect 1857 1192 1887 1218
rect 1953 1196 1983 1218
rect 1743 1146 1759 1180
rect 1793 1146 1809 1180
rect 1743 1130 1809 1146
rect 1935 1180 2001 1196
rect 2049 1192 2079 1218
rect 2145 1196 2175 1218
rect 1935 1146 1951 1180
rect 1985 1146 2001 1180
rect 1935 1130 2001 1146
rect 2127 1180 2193 1196
rect 2241 1192 2271 1218
rect 2337 1196 2367 1218
rect 2127 1146 2143 1180
rect 2177 1146 2193 1180
rect 2127 1130 2193 1146
rect 2319 1180 2385 1196
rect 2433 1192 2463 1218
rect 2529 1196 2559 1218
rect 2319 1146 2335 1180
rect 2369 1146 2385 1180
rect 2319 1130 2385 1146
rect 2511 1180 2577 1196
rect 2625 1192 2655 1218
rect 2721 1196 2751 1218
rect 2511 1146 2527 1180
rect 2561 1146 2577 1180
rect 2511 1130 2577 1146
rect 2703 1180 2769 1196
rect 2817 1192 2847 1218
rect 2703 1146 2719 1180
rect 2753 1146 2769 1180
rect 2703 1130 2769 1146
rect -2865 1072 -2799 1088
rect -2865 1038 -2849 1072
rect -2815 1038 -2799 1072
rect -2865 1022 -2799 1038
rect -2673 1072 -2607 1088
rect -2673 1038 -2657 1072
rect -2623 1038 -2607 1072
rect -2847 1000 -2817 1022
rect -2751 1000 -2721 1026
rect -2673 1022 -2607 1038
rect -2481 1072 -2415 1088
rect -2481 1038 -2465 1072
rect -2431 1038 -2415 1072
rect -2655 1000 -2625 1022
rect -2559 1000 -2529 1026
rect -2481 1022 -2415 1038
rect -2289 1072 -2223 1088
rect -2289 1038 -2273 1072
rect -2239 1038 -2223 1072
rect -2463 1000 -2433 1022
rect -2367 1000 -2337 1026
rect -2289 1022 -2223 1038
rect -2097 1072 -2031 1088
rect -2097 1038 -2081 1072
rect -2047 1038 -2031 1072
rect -2271 1000 -2241 1022
rect -2175 1000 -2145 1026
rect -2097 1022 -2031 1038
rect -1905 1072 -1839 1088
rect -1905 1038 -1889 1072
rect -1855 1038 -1839 1072
rect -2079 1000 -2049 1022
rect -1983 1000 -1953 1026
rect -1905 1022 -1839 1038
rect -1713 1072 -1647 1088
rect -1713 1038 -1697 1072
rect -1663 1038 -1647 1072
rect -1887 1000 -1857 1022
rect -1791 1000 -1761 1026
rect -1713 1022 -1647 1038
rect -1521 1072 -1455 1088
rect -1521 1038 -1505 1072
rect -1471 1038 -1455 1072
rect -1695 1000 -1665 1022
rect -1599 1000 -1569 1026
rect -1521 1022 -1455 1038
rect -1329 1072 -1263 1088
rect -1329 1038 -1313 1072
rect -1279 1038 -1263 1072
rect -1503 1000 -1473 1022
rect -1407 1000 -1377 1026
rect -1329 1022 -1263 1038
rect -1137 1072 -1071 1088
rect -1137 1038 -1121 1072
rect -1087 1038 -1071 1072
rect -1311 1000 -1281 1022
rect -1215 1000 -1185 1026
rect -1137 1022 -1071 1038
rect -945 1072 -879 1088
rect -945 1038 -929 1072
rect -895 1038 -879 1072
rect -1119 1000 -1089 1022
rect -1023 1000 -993 1026
rect -945 1022 -879 1038
rect -753 1072 -687 1088
rect -753 1038 -737 1072
rect -703 1038 -687 1072
rect -927 1000 -897 1022
rect -831 1000 -801 1026
rect -753 1022 -687 1038
rect -561 1072 -495 1088
rect -561 1038 -545 1072
rect -511 1038 -495 1072
rect -735 1000 -705 1022
rect -639 1000 -609 1026
rect -561 1022 -495 1038
rect -369 1072 -303 1088
rect -369 1038 -353 1072
rect -319 1038 -303 1072
rect -543 1000 -513 1022
rect -447 1000 -417 1026
rect -369 1022 -303 1038
rect -177 1072 -111 1088
rect -177 1038 -161 1072
rect -127 1038 -111 1072
rect -351 1000 -321 1022
rect -255 1000 -225 1026
rect -177 1022 -111 1038
rect 15 1072 81 1088
rect 15 1038 31 1072
rect 65 1038 81 1072
rect -159 1000 -129 1022
rect -63 1000 -33 1026
rect 15 1022 81 1038
rect 207 1072 273 1088
rect 207 1038 223 1072
rect 257 1038 273 1072
rect 33 1000 63 1022
rect 129 1000 159 1026
rect 207 1022 273 1038
rect 399 1072 465 1088
rect 399 1038 415 1072
rect 449 1038 465 1072
rect 225 1000 255 1022
rect 321 1000 351 1026
rect 399 1022 465 1038
rect 591 1072 657 1088
rect 591 1038 607 1072
rect 641 1038 657 1072
rect 417 1000 447 1022
rect 513 1000 543 1026
rect 591 1022 657 1038
rect 783 1072 849 1088
rect 783 1038 799 1072
rect 833 1038 849 1072
rect 609 1000 639 1022
rect 705 1000 735 1026
rect 783 1022 849 1038
rect 975 1072 1041 1088
rect 975 1038 991 1072
rect 1025 1038 1041 1072
rect 801 1000 831 1022
rect 897 1000 927 1026
rect 975 1022 1041 1038
rect 1167 1072 1233 1088
rect 1167 1038 1183 1072
rect 1217 1038 1233 1072
rect 993 1000 1023 1022
rect 1089 1000 1119 1026
rect 1167 1022 1233 1038
rect 1359 1072 1425 1088
rect 1359 1038 1375 1072
rect 1409 1038 1425 1072
rect 1185 1000 1215 1022
rect 1281 1000 1311 1026
rect 1359 1022 1425 1038
rect 1551 1072 1617 1088
rect 1551 1038 1567 1072
rect 1601 1038 1617 1072
rect 1377 1000 1407 1022
rect 1473 1000 1503 1026
rect 1551 1022 1617 1038
rect 1743 1072 1809 1088
rect 1743 1038 1759 1072
rect 1793 1038 1809 1072
rect 1569 1000 1599 1022
rect 1665 1000 1695 1026
rect 1743 1022 1809 1038
rect 1935 1072 2001 1088
rect 1935 1038 1951 1072
rect 1985 1038 2001 1072
rect 1761 1000 1791 1022
rect 1857 1000 1887 1026
rect 1935 1022 2001 1038
rect 2127 1072 2193 1088
rect 2127 1038 2143 1072
rect 2177 1038 2193 1072
rect 1953 1000 1983 1022
rect 2049 1000 2079 1026
rect 2127 1022 2193 1038
rect 2319 1072 2385 1088
rect 2319 1038 2335 1072
rect 2369 1038 2385 1072
rect 2145 1000 2175 1022
rect 2241 1000 2271 1026
rect 2319 1022 2385 1038
rect 2511 1072 2577 1088
rect 2511 1038 2527 1072
rect 2561 1038 2577 1072
rect 2337 1000 2367 1022
rect 2433 1000 2463 1026
rect 2511 1022 2577 1038
rect 2703 1072 2769 1088
rect 2703 1038 2719 1072
rect 2753 1038 2769 1072
rect 2529 1000 2559 1022
rect 2625 1000 2655 1026
rect 2703 1022 2769 1038
rect 2721 1000 2751 1022
rect 2817 1000 2847 1026
rect -2847 -1026 -2817 -1000
rect -2751 -1022 -2721 -1000
rect -2769 -1038 -2703 -1022
rect -2655 -1026 -2625 -1000
rect -2559 -1022 -2529 -1000
rect -2769 -1072 -2753 -1038
rect -2719 -1072 -2703 -1038
rect -2769 -1088 -2703 -1072
rect -2577 -1038 -2511 -1022
rect -2463 -1026 -2433 -1000
rect -2367 -1022 -2337 -1000
rect -2577 -1072 -2561 -1038
rect -2527 -1072 -2511 -1038
rect -2577 -1088 -2511 -1072
rect -2385 -1038 -2319 -1022
rect -2271 -1026 -2241 -1000
rect -2175 -1022 -2145 -1000
rect -2385 -1072 -2369 -1038
rect -2335 -1072 -2319 -1038
rect -2385 -1088 -2319 -1072
rect -2193 -1038 -2127 -1022
rect -2079 -1026 -2049 -1000
rect -1983 -1022 -1953 -1000
rect -2193 -1072 -2177 -1038
rect -2143 -1072 -2127 -1038
rect -2193 -1088 -2127 -1072
rect -2001 -1038 -1935 -1022
rect -1887 -1026 -1857 -1000
rect -1791 -1022 -1761 -1000
rect -2001 -1072 -1985 -1038
rect -1951 -1072 -1935 -1038
rect -2001 -1088 -1935 -1072
rect -1809 -1038 -1743 -1022
rect -1695 -1026 -1665 -1000
rect -1599 -1022 -1569 -1000
rect -1809 -1072 -1793 -1038
rect -1759 -1072 -1743 -1038
rect -1809 -1088 -1743 -1072
rect -1617 -1038 -1551 -1022
rect -1503 -1026 -1473 -1000
rect -1407 -1022 -1377 -1000
rect -1617 -1072 -1601 -1038
rect -1567 -1072 -1551 -1038
rect -1617 -1088 -1551 -1072
rect -1425 -1038 -1359 -1022
rect -1311 -1026 -1281 -1000
rect -1215 -1022 -1185 -1000
rect -1425 -1072 -1409 -1038
rect -1375 -1072 -1359 -1038
rect -1425 -1088 -1359 -1072
rect -1233 -1038 -1167 -1022
rect -1119 -1026 -1089 -1000
rect -1023 -1022 -993 -1000
rect -1233 -1072 -1217 -1038
rect -1183 -1072 -1167 -1038
rect -1233 -1088 -1167 -1072
rect -1041 -1038 -975 -1022
rect -927 -1026 -897 -1000
rect -831 -1022 -801 -1000
rect -1041 -1072 -1025 -1038
rect -991 -1072 -975 -1038
rect -1041 -1088 -975 -1072
rect -849 -1038 -783 -1022
rect -735 -1026 -705 -1000
rect -639 -1022 -609 -1000
rect -849 -1072 -833 -1038
rect -799 -1072 -783 -1038
rect -849 -1088 -783 -1072
rect -657 -1038 -591 -1022
rect -543 -1026 -513 -1000
rect -447 -1022 -417 -1000
rect -657 -1072 -641 -1038
rect -607 -1072 -591 -1038
rect -657 -1088 -591 -1072
rect -465 -1038 -399 -1022
rect -351 -1026 -321 -1000
rect -255 -1022 -225 -1000
rect -465 -1072 -449 -1038
rect -415 -1072 -399 -1038
rect -465 -1088 -399 -1072
rect -273 -1038 -207 -1022
rect -159 -1026 -129 -1000
rect -63 -1022 -33 -1000
rect -273 -1072 -257 -1038
rect -223 -1072 -207 -1038
rect -273 -1088 -207 -1072
rect -81 -1038 -15 -1022
rect 33 -1026 63 -1000
rect 129 -1022 159 -1000
rect -81 -1072 -65 -1038
rect -31 -1072 -15 -1038
rect -81 -1088 -15 -1072
rect 111 -1038 177 -1022
rect 225 -1026 255 -1000
rect 321 -1022 351 -1000
rect 111 -1072 127 -1038
rect 161 -1072 177 -1038
rect 111 -1088 177 -1072
rect 303 -1038 369 -1022
rect 417 -1026 447 -1000
rect 513 -1022 543 -1000
rect 303 -1072 319 -1038
rect 353 -1072 369 -1038
rect 303 -1088 369 -1072
rect 495 -1038 561 -1022
rect 609 -1026 639 -1000
rect 705 -1022 735 -1000
rect 495 -1072 511 -1038
rect 545 -1072 561 -1038
rect 495 -1088 561 -1072
rect 687 -1038 753 -1022
rect 801 -1026 831 -1000
rect 897 -1022 927 -1000
rect 687 -1072 703 -1038
rect 737 -1072 753 -1038
rect 687 -1088 753 -1072
rect 879 -1038 945 -1022
rect 993 -1026 1023 -1000
rect 1089 -1022 1119 -1000
rect 879 -1072 895 -1038
rect 929 -1072 945 -1038
rect 879 -1088 945 -1072
rect 1071 -1038 1137 -1022
rect 1185 -1026 1215 -1000
rect 1281 -1022 1311 -1000
rect 1071 -1072 1087 -1038
rect 1121 -1072 1137 -1038
rect 1071 -1088 1137 -1072
rect 1263 -1038 1329 -1022
rect 1377 -1026 1407 -1000
rect 1473 -1022 1503 -1000
rect 1263 -1072 1279 -1038
rect 1313 -1072 1329 -1038
rect 1263 -1088 1329 -1072
rect 1455 -1038 1521 -1022
rect 1569 -1026 1599 -1000
rect 1665 -1022 1695 -1000
rect 1455 -1072 1471 -1038
rect 1505 -1072 1521 -1038
rect 1455 -1088 1521 -1072
rect 1647 -1038 1713 -1022
rect 1761 -1026 1791 -1000
rect 1857 -1022 1887 -1000
rect 1647 -1072 1663 -1038
rect 1697 -1072 1713 -1038
rect 1647 -1088 1713 -1072
rect 1839 -1038 1905 -1022
rect 1953 -1026 1983 -1000
rect 2049 -1022 2079 -1000
rect 1839 -1072 1855 -1038
rect 1889 -1072 1905 -1038
rect 1839 -1088 1905 -1072
rect 2031 -1038 2097 -1022
rect 2145 -1026 2175 -1000
rect 2241 -1022 2271 -1000
rect 2031 -1072 2047 -1038
rect 2081 -1072 2097 -1038
rect 2031 -1088 2097 -1072
rect 2223 -1038 2289 -1022
rect 2337 -1026 2367 -1000
rect 2433 -1022 2463 -1000
rect 2223 -1072 2239 -1038
rect 2273 -1072 2289 -1038
rect 2223 -1088 2289 -1072
rect 2415 -1038 2481 -1022
rect 2529 -1026 2559 -1000
rect 2625 -1022 2655 -1000
rect 2415 -1072 2431 -1038
rect 2465 -1072 2481 -1038
rect 2415 -1088 2481 -1072
rect 2607 -1038 2673 -1022
rect 2721 -1026 2751 -1000
rect 2817 -1022 2847 -1000
rect 2607 -1072 2623 -1038
rect 2657 -1072 2673 -1038
rect 2607 -1088 2673 -1072
rect 2799 -1038 2865 -1022
rect 2799 -1072 2815 -1038
rect 2849 -1072 2865 -1038
rect 2799 -1088 2865 -1072
rect -2769 -1146 -2703 -1130
rect -2769 -1180 -2753 -1146
rect -2719 -1180 -2703 -1146
rect -2847 -1218 -2817 -1192
rect -2769 -1196 -2703 -1180
rect -2577 -1146 -2511 -1130
rect -2577 -1180 -2561 -1146
rect -2527 -1180 -2511 -1146
rect -2751 -1218 -2721 -1196
rect -2655 -1218 -2625 -1192
rect -2577 -1196 -2511 -1180
rect -2385 -1146 -2319 -1130
rect -2385 -1180 -2369 -1146
rect -2335 -1180 -2319 -1146
rect -2559 -1218 -2529 -1196
rect -2463 -1218 -2433 -1192
rect -2385 -1196 -2319 -1180
rect -2193 -1146 -2127 -1130
rect -2193 -1180 -2177 -1146
rect -2143 -1180 -2127 -1146
rect -2367 -1218 -2337 -1196
rect -2271 -1218 -2241 -1192
rect -2193 -1196 -2127 -1180
rect -2001 -1146 -1935 -1130
rect -2001 -1180 -1985 -1146
rect -1951 -1180 -1935 -1146
rect -2175 -1218 -2145 -1196
rect -2079 -1218 -2049 -1192
rect -2001 -1196 -1935 -1180
rect -1809 -1146 -1743 -1130
rect -1809 -1180 -1793 -1146
rect -1759 -1180 -1743 -1146
rect -1983 -1218 -1953 -1196
rect -1887 -1218 -1857 -1192
rect -1809 -1196 -1743 -1180
rect -1617 -1146 -1551 -1130
rect -1617 -1180 -1601 -1146
rect -1567 -1180 -1551 -1146
rect -1791 -1218 -1761 -1196
rect -1695 -1218 -1665 -1192
rect -1617 -1196 -1551 -1180
rect -1425 -1146 -1359 -1130
rect -1425 -1180 -1409 -1146
rect -1375 -1180 -1359 -1146
rect -1599 -1218 -1569 -1196
rect -1503 -1218 -1473 -1192
rect -1425 -1196 -1359 -1180
rect -1233 -1146 -1167 -1130
rect -1233 -1180 -1217 -1146
rect -1183 -1180 -1167 -1146
rect -1407 -1218 -1377 -1196
rect -1311 -1218 -1281 -1192
rect -1233 -1196 -1167 -1180
rect -1041 -1146 -975 -1130
rect -1041 -1180 -1025 -1146
rect -991 -1180 -975 -1146
rect -1215 -1218 -1185 -1196
rect -1119 -1218 -1089 -1192
rect -1041 -1196 -975 -1180
rect -849 -1146 -783 -1130
rect -849 -1180 -833 -1146
rect -799 -1180 -783 -1146
rect -1023 -1218 -993 -1196
rect -927 -1218 -897 -1192
rect -849 -1196 -783 -1180
rect -657 -1146 -591 -1130
rect -657 -1180 -641 -1146
rect -607 -1180 -591 -1146
rect -831 -1218 -801 -1196
rect -735 -1218 -705 -1192
rect -657 -1196 -591 -1180
rect -465 -1146 -399 -1130
rect -465 -1180 -449 -1146
rect -415 -1180 -399 -1146
rect -639 -1218 -609 -1196
rect -543 -1218 -513 -1192
rect -465 -1196 -399 -1180
rect -273 -1146 -207 -1130
rect -273 -1180 -257 -1146
rect -223 -1180 -207 -1146
rect -447 -1218 -417 -1196
rect -351 -1218 -321 -1192
rect -273 -1196 -207 -1180
rect -81 -1146 -15 -1130
rect -81 -1180 -65 -1146
rect -31 -1180 -15 -1146
rect -255 -1218 -225 -1196
rect -159 -1218 -129 -1192
rect -81 -1196 -15 -1180
rect 111 -1146 177 -1130
rect 111 -1180 127 -1146
rect 161 -1180 177 -1146
rect -63 -1218 -33 -1196
rect 33 -1218 63 -1192
rect 111 -1196 177 -1180
rect 303 -1146 369 -1130
rect 303 -1180 319 -1146
rect 353 -1180 369 -1146
rect 129 -1218 159 -1196
rect 225 -1218 255 -1192
rect 303 -1196 369 -1180
rect 495 -1146 561 -1130
rect 495 -1180 511 -1146
rect 545 -1180 561 -1146
rect 321 -1218 351 -1196
rect 417 -1218 447 -1192
rect 495 -1196 561 -1180
rect 687 -1146 753 -1130
rect 687 -1180 703 -1146
rect 737 -1180 753 -1146
rect 513 -1218 543 -1196
rect 609 -1218 639 -1192
rect 687 -1196 753 -1180
rect 879 -1146 945 -1130
rect 879 -1180 895 -1146
rect 929 -1180 945 -1146
rect 705 -1218 735 -1196
rect 801 -1218 831 -1192
rect 879 -1196 945 -1180
rect 1071 -1146 1137 -1130
rect 1071 -1180 1087 -1146
rect 1121 -1180 1137 -1146
rect 897 -1218 927 -1196
rect 993 -1218 1023 -1192
rect 1071 -1196 1137 -1180
rect 1263 -1146 1329 -1130
rect 1263 -1180 1279 -1146
rect 1313 -1180 1329 -1146
rect 1089 -1218 1119 -1196
rect 1185 -1218 1215 -1192
rect 1263 -1196 1329 -1180
rect 1455 -1146 1521 -1130
rect 1455 -1180 1471 -1146
rect 1505 -1180 1521 -1146
rect 1281 -1218 1311 -1196
rect 1377 -1218 1407 -1192
rect 1455 -1196 1521 -1180
rect 1647 -1146 1713 -1130
rect 1647 -1180 1663 -1146
rect 1697 -1180 1713 -1146
rect 1473 -1218 1503 -1196
rect 1569 -1218 1599 -1192
rect 1647 -1196 1713 -1180
rect 1839 -1146 1905 -1130
rect 1839 -1180 1855 -1146
rect 1889 -1180 1905 -1146
rect 1665 -1218 1695 -1196
rect 1761 -1218 1791 -1192
rect 1839 -1196 1905 -1180
rect 2031 -1146 2097 -1130
rect 2031 -1180 2047 -1146
rect 2081 -1180 2097 -1146
rect 1857 -1218 1887 -1196
rect 1953 -1218 1983 -1192
rect 2031 -1196 2097 -1180
rect 2223 -1146 2289 -1130
rect 2223 -1180 2239 -1146
rect 2273 -1180 2289 -1146
rect 2049 -1218 2079 -1196
rect 2145 -1218 2175 -1192
rect 2223 -1196 2289 -1180
rect 2415 -1146 2481 -1130
rect 2415 -1180 2431 -1146
rect 2465 -1180 2481 -1146
rect 2241 -1218 2271 -1196
rect 2337 -1218 2367 -1192
rect 2415 -1196 2481 -1180
rect 2607 -1146 2673 -1130
rect 2607 -1180 2623 -1146
rect 2657 -1180 2673 -1146
rect 2433 -1218 2463 -1196
rect 2529 -1218 2559 -1192
rect 2607 -1196 2673 -1180
rect 2799 -1146 2865 -1130
rect 2799 -1180 2815 -1146
rect 2849 -1180 2865 -1146
rect 2625 -1218 2655 -1196
rect 2721 -1218 2751 -1192
rect 2799 -1196 2865 -1180
rect 2817 -1218 2847 -1196
rect -2847 -3240 -2817 -3218
rect -2865 -3256 -2799 -3240
rect -2751 -3244 -2721 -3218
rect -2655 -3240 -2625 -3218
rect -2865 -3290 -2849 -3256
rect -2815 -3290 -2799 -3256
rect -2865 -3306 -2799 -3290
rect -2673 -3256 -2607 -3240
rect -2559 -3244 -2529 -3218
rect -2463 -3240 -2433 -3218
rect -2673 -3290 -2657 -3256
rect -2623 -3290 -2607 -3256
rect -2673 -3306 -2607 -3290
rect -2481 -3256 -2415 -3240
rect -2367 -3244 -2337 -3218
rect -2271 -3240 -2241 -3218
rect -2481 -3290 -2465 -3256
rect -2431 -3290 -2415 -3256
rect -2481 -3306 -2415 -3290
rect -2289 -3256 -2223 -3240
rect -2175 -3244 -2145 -3218
rect -2079 -3240 -2049 -3218
rect -2289 -3290 -2273 -3256
rect -2239 -3290 -2223 -3256
rect -2289 -3306 -2223 -3290
rect -2097 -3256 -2031 -3240
rect -1983 -3244 -1953 -3218
rect -1887 -3240 -1857 -3218
rect -2097 -3290 -2081 -3256
rect -2047 -3290 -2031 -3256
rect -2097 -3306 -2031 -3290
rect -1905 -3256 -1839 -3240
rect -1791 -3244 -1761 -3218
rect -1695 -3240 -1665 -3218
rect -1905 -3290 -1889 -3256
rect -1855 -3290 -1839 -3256
rect -1905 -3306 -1839 -3290
rect -1713 -3256 -1647 -3240
rect -1599 -3244 -1569 -3218
rect -1503 -3240 -1473 -3218
rect -1713 -3290 -1697 -3256
rect -1663 -3290 -1647 -3256
rect -1713 -3306 -1647 -3290
rect -1521 -3256 -1455 -3240
rect -1407 -3244 -1377 -3218
rect -1311 -3240 -1281 -3218
rect -1521 -3290 -1505 -3256
rect -1471 -3290 -1455 -3256
rect -1521 -3306 -1455 -3290
rect -1329 -3256 -1263 -3240
rect -1215 -3244 -1185 -3218
rect -1119 -3240 -1089 -3218
rect -1329 -3290 -1313 -3256
rect -1279 -3290 -1263 -3256
rect -1329 -3306 -1263 -3290
rect -1137 -3256 -1071 -3240
rect -1023 -3244 -993 -3218
rect -927 -3240 -897 -3218
rect -1137 -3290 -1121 -3256
rect -1087 -3290 -1071 -3256
rect -1137 -3306 -1071 -3290
rect -945 -3256 -879 -3240
rect -831 -3244 -801 -3218
rect -735 -3240 -705 -3218
rect -945 -3290 -929 -3256
rect -895 -3290 -879 -3256
rect -945 -3306 -879 -3290
rect -753 -3256 -687 -3240
rect -639 -3244 -609 -3218
rect -543 -3240 -513 -3218
rect -753 -3290 -737 -3256
rect -703 -3290 -687 -3256
rect -753 -3306 -687 -3290
rect -561 -3256 -495 -3240
rect -447 -3244 -417 -3218
rect -351 -3240 -321 -3218
rect -561 -3290 -545 -3256
rect -511 -3290 -495 -3256
rect -561 -3306 -495 -3290
rect -369 -3256 -303 -3240
rect -255 -3244 -225 -3218
rect -159 -3240 -129 -3218
rect -369 -3290 -353 -3256
rect -319 -3290 -303 -3256
rect -369 -3306 -303 -3290
rect -177 -3256 -111 -3240
rect -63 -3244 -33 -3218
rect 33 -3240 63 -3218
rect -177 -3290 -161 -3256
rect -127 -3290 -111 -3256
rect -177 -3306 -111 -3290
rect 15 -3256 81 -3240
rect 129 -3244 159 -3218
rect 225 -3240 255 -3218
rect 15 -3290 31 -3256
rect 65 -3290 81 -3256
rect 15 -3306 81 -3290
rect 207 -3256 273 -3240
rect 321 -3244 351 -3218
rect 417 -3240 447 -3218
rect 207 -3290 223 -3256
rect 257 -3290 273 -3256
rect 207 -3306 273 -3290
rect 399 -3256 465 -3240
rect 513 -3244 543 -3218
rect 609 -3240 639 -3218
rect 399 -3290 415 -3256
rect 449 -3290 465 -3256
rect 399 -3306 465 -3290
rect 591 -3256 657 -3240
rect 705 -3244 735 -3218
rect 801 -3240 831 -3218
rect 591 -3290 607 -3256
rect 641 -3290 657 -3256
rect 591 -3306 657 -3290
rect 783 -3256 849 -3240
rect 897 -3244 927 -3218
rect 993 -3240 1023 -3218
rect 783 -3290 799 -3256
rect 833 -3290 849 -3256
rect 783 -3306 849 -3290
rect 975 -3256 1041 -3240
rect 1089 -3244 1119 -3218
rect 1185 -3240 1215 -3218
rect 975 -3290 991 -3256
rect 1025 -3290 1041 -3256
rect 975 -3306 1041 -3290
rect 1167 -3256 1233 -3240
rect 1281 -3244 1311 -3218
rect 1377 -3240 1407 -3218
rect 1167 -3290 1183 -3256
rect 1217 -3290 1233 -3256
rect 1167 -3306 1233 -3290
rect 1359 -3256 1425 -3240
rect 1473 -3244 1503 -3218
rect 1569 -3240 1599 -3218
rect 1359 -3290 1375 -3256
rect 1409 -3290 1425 -3256
rect 1359 -3306 1425 -3290
rect 1551 -3256 1617 -3240
rect 1665 -3244 1695 -3218
rect 1761 -3240 1791 -3218
rect 1551 -3290 1567 -3256
rect 1601 -3290 1617 -3256
rect 1551 -3306 1617 -3290
rect 1743 -3256 1809 -3240
rect 1857 -3244 1887 -3218
rect 1953 -3240 1983 -3218
rect 1743 -3290 1759 -3256
rect 1793 -3290 1809 -3256
rect 1743 -3306 1809 -3290
rect 1935 -3256 2001 -3240
rect 2049 -3244 2079 -3218
rect 2145 -3240 2175 -3218
rect 1935 -3290 1951 -3256
rect 1985 -3290 2001 -3256
rect 1935 -3306 2001 -3290
rect 2127 -3256 2193 -3240
rect 2241 -3244 2271 -3218
rect 2337 -3240 2367 -3218
rect 2127 -3290 2143 -3256
rect 2177 -3290 2193 -3256
rect 2127 -3306 2193 -3290
rect 2319 -3256 2385 -3240
rect 2433 -3244 2463 -3218
rect 2529 -3240 2559 -3218
rect 2319 -3290 2335 -3256
rect 2369 -3290 2385 -3256
rect 2319 -3306 2385 -3290
rect 2511 -3256 2577 -3240
rect 2625 -3244 2655 -3218
rect 2721 -3240 2751 -3218
rect 2511 -3290 2527 -3256
rect 2561 -3290 2577 -3256
rect 2511 -3306 2577 -3290
rect 2703 -3256 2769 -3240
rect 2817 -3244 2847 -3218
rect 2703 -3290 2719 -3256
rect 2753 -3290 2769 -3256
rect 2703 -3306 2769 -3290
<< polycont >>
rect -2753 3256 -2719 3290
rect -2561 3256 -2527 3290
rect -2369 3256 -2335 3290
rect -2177 3256 -2143 3290
rect -1985 3256 -1951 3290
rect -1793 3256 -1759 3290
rect -1601 3256 -1567 3290
rect -1409 3256 -1375 3290
rect -1217 3256 -1183 3290
rect -1025 3256 -991 3290
rect -833 3256 -799 3290
rect -641 3256 -607 3290
rect -449 3256 -415 3290
rect -257 3256 -223 3290
rect -65 3256 -31 3290
rect 127 3256 161 3290
rect 319 3256 353 3290
rect 511 3256 545 3290
rect 703 3256 737 3290
rect 895 3256 929 3290
rect 1087 3256 1121 3290
rect 1279 3256 1313 3290
rect 1471 3256 1505 3290
rect 1663 3256 1697 3290
rect 1855 3256 1889 3290
rect 2047 3256 2081 3290
rect 2239 3256 2273 3290
rect 2431 3256 2465 3290
rect 2623 3256 2657 3290
rect 2815 3256 2849 3290
rect -2849 1146 -2815 1180
rect -2657 1146 -2623 1180
rect -2465 1146 -2431 1180
rect -2273 1146 -2239 1180
rect -2081 1146 -2047 1180
rect -1889 1146 -1855 1180
rect -1697 1146 -1663 1180
rect -1505 1146 -1471 1180
rect -1313 1146 -1279 1180
rect -1121 1146 -1087 1180
rect -929 1146 -895 1180
rect -737 1146 -703 1180
rect -545 1146 -511 1180
rect -353 1146 -319 1180
rect -161 1146 -127 1180
rect 31 1146 65 1180
rect 223 1146 257 1180
rect 415 1146 449 1180
rect 607 1146 641 1180
rect 799 1146 833 1180
rect 991 1146 1025 1180
rect 1183 1146 1217 1180
rect 1375 1146 1409 1180
rect 1567 1146 1601 1180
rect 1759 1146 1793 1180
rect 1951 1146 1985 1180
rect 2143 1146 2177 1180
rect 2335 1146 2369 1180
rect 2527 1146 2561 1180
rect 2719 1146 2753 1180
rect -2849 1038 -2815 1072
rect -2657 1038 -2623 1072
rect -2465 1038 -2431 1072
rect -2273 1038 -2239 1072
rect -2081 1038 -2047 1072
rect -1889 1038 -1855 1072
rect -1697 1038 -1663 1072
rect -1505 1038 -1471 1072
rect -1313 1038 -1279 1072
rect -1121 1038 -1087 1072
rect -929 1038 -895 1072
rect -737 1038 -703 1072
rect -545 1038 -511 1072
rect -353 1038 -319 1072
rect -161 1038 -127 1072
rect 31 1038 65 1072
rect 223 1038 257 1072
rect 415 1038 449 1072
rect 607 1038 641 1072
rect 799 1038 833 1072
rect 991 1038 1025 1072
rect 1183 1038 1217 1072
rect 1375 1038 1409 1072
rect 1567 1038 1601 1072
rect 1759 1038 1793 1072
rect 1951 1038 1985 1072
rect 2143 1038 2177 1072
rect 2335 1038 2369 1072
rect 2527 1038 2561 1072
rect 2719 1038 2753 1072
rect -2753 -1072 -2719 -1038
rect -2561 -1072 -2527 -1038
rect -2369 -1072 -2335 -1038
rect -2177 -1072 -2143 -1038
rect -1985 -1072 -1951 -1038
rect -1793 -1072 -1759 -1038
rect -1601 -1072 -1567 -1038
rect -1409 -1072 -1375 -1038
rect -1217 -1072 -1183 -1038
rect -1025 -1072 -991 -1038
rect -833 -1072 -799 -1038
rect -641 -1072 -607 -1038
rect -449 -1072 -415 -1038
rect -257 -1072 -223 -1038
rect -65 -1072 -31 -1038
rect 127 -1072 161 -1038
rect 319 -1072 353 -1038
rect 511 -1072 545 -1038
rect 703 -1072 737 -1038
rect 895 -1072 929 -1038
rect 1087 -1072 1121 -1038
rect 1279 -1072 1313 -1038
rect 1471 -1072 1505 -1038
rect 1663 -1072 1697 -1038
rect 1855 -1072 1889 -1038
rect 2047 -1072 2081 -1038
rect 2239 -1072 2273 -1038
rect 2431 -1072 2465 -1038
rect 2623 -1072 2657 -1038
rect 2815 -1072 2849 -1038
rect -2753 -1180 -2719 -1146
rect -2561 -1180 -2527 -1146
rect -2369 -1180 -2335 -1146
rect -2177 -1180 -2143 -1146
rect -1985 -1180 -1951 -1146
rect -1793 -1180 -1759 -1146
rect -1601 -1180 -1567 -1146
rect -1409 -1180 -1375 -1146
rect -1217 -1180 -1183 -1146
rect -1025 -1180 -991 -1146
rect -833 -1180 -799 -1146
rect -641 -1180 -607 -1146
rect -449 -1180 -415 -1146
rect -257 -1180 -223 -1146
rect -65 -1180 -31 -1146
rect 127 -1180 161 -1146
rect 319 -1180 353 -1146
rect 511 -1180 545 -1146
rect 703 -1180 737 -1146
rect 895 -1180 929 -1146
rect 1087 -1180 1121 -1146
rect 1279 -1180 1313 -1146
rect 1471 -1180 1505 -1146
rect 1663 -1180 1697 -1146
rect 1855 -1180 1889 -1146
rect 2047 -1180 2081 -1146
rect 2239 -1180 2273 -1146
rect 2431 -1180 2465 -1146
rect 2623 -1180 2657 -1146
rect 2815 -1180 2849 -1146
rect -2849 -3290 -2815 -3256
rect -2657 -3290 -2623 -3256
rect -2465 -3290 -2431 -3256
rect -2273 -3290 -2239 -3256
rect -2081 -3290 -2047 -3256
rect -1889 -3290 -1855 -3256
rect -1697 -3290 -1663 -3256
rect -1505 -3290 -1471 -3256
rect -1313 -3290 -1279 -3256
rect -1121 -3290 -1087 -3256
rect -929 -3290 -895 -3256
rect -737 -3290 -703 -3256
rect -545 -3290 -511 -3256
rect -353 -3290 -319 -3256
rect -161 -3290 -127 -3256
rect 31 -3290 65 -3256
rect 223 -3290 257 -3256
rect 415 -3290 449 -3256
rect 607 -3290 641 -3256
rect 799 -3290 833 -3256
rect 991 -3290 1025 -3256
rect 1183 -3290 1217 -3256
rect 1375 -3290 1409 -3256
rect 1567 -3290 1601 -3256
rect 1759 -3290 1793 -3256
rect 1951 -3290 1985 -3256
rect 2143 -3290 2177 -3256
rect 2335 -3290 2369 -3256
rect 2527 -3290 2561 -3256
rect 2719 -3290 2753 -3256
<< locali >>
rect -2769 3256 -2753 3290
rect -2719 3256 -2703 3290
rect -2577 3256 -2561 3290
rect -2527 3256 -2511 3290
rect -2385 3256 -2369 3290
rect -2335 3256 -2319 3290
rect -2193 3256 -2177 3290
rect -2143 3256 -2127 3290
rect -2001 3256 -1985 3290
rect -1951 3256 -1935 3290
rect -1809 3256 -1793 3290
rect -1759 3256 -1743 3290
rect -1617 3256 -1601 3290
rect -1567 3256 -1551 3290
rect -1425 3256 -1409 3290
rect -1375 3256 -1359 3290
rect -1233 3256 -1217 3290
rect -1183 3256 -1167 3290
rect -1041 3256 -1025 3290
rect -991 3256 -975 3290
rect -849 3256 -833 3290
rect -799 3256 -783 3290
rect -657 3256 -641 3290
rect -607 3256 -591 3290
rect -465 3256 -449 3290
rect -415 3256 -399 3290
rect -273 3256 -257 3290
rect -223 3256 -207 3290
rect -81 3256 -65 3290
rect -31 3256 -15 3290
rect 111 3256 127 3290
rect 161 3256 177 3290
rect 303 3256 319 3290
rect 353 3256 369 3290
rect 495 3256 511 3290
rect 545 3256 561 3290
rect 687 3256 703 3290
rect 737 3256 753 3290
rect 879 3256 895 3290
rect 929 3256 945 3290
rect 1071 3256 1087 3290
rect 1121 3256 1137 3290
rect 1263 3256 1279 3290
rect 1313 3256 1329 3290
rect 1455 3256 1471 3290
rect 1505 3256 1521 3290
rect 1647 3256 1663 3290
rect 1697 3256 1713 3290
rect 1839 3256 1855 3290
rect 1889 3256 1905 3290
rect 2031 3256 2047 3290
rect 2081 3256 2097 3290
rect 2223 3256 2239 3290
rect 2273 3256 2289 3290
rect 2415 3256 2431 3290
rect 2465 3256 2481 3290
rect 2607 3256 2623 3290
rect 2657 3256 2673 3290
rect 2799 3256 2815 3290
rect 2849 3256 2865 3290
rect -2897 3206 -2863 3222
rect -2897 1214 -2863 1230
rect -2801 3206 -2767 3222
rect -2801 1214 -2767 1230
rect -2705 3206 -2671 3222
rect -2705 1214 -2671 1230
rect -2609 3206 -2575 3222
rect -2609 1214 -2575 1230
rect -2513 3206 -2479 3222
rect -2513 1214 -2479 1230
rect -2417 3206 -2383 3222
rect -2417 1214 -2383 1230
rect -2321 3206 -2287 3222
rect -2321 1214 -2287 1230
rect -2225 3206 -2191 3222
rect -2225 1214 -2191 1230
rect -2129 3206 -2095 3222
rect -2129 1214 -2095 1230
rect -2033 3206 -1999 3222
rect -2033 1214 -1999 1230
rect -1937 3206 -1903 3222
rect -1937 1214 -1903 1230
rect -1841 3206 -1807 3222
rect -1841 1214 -1807 1230
rect -1745 3206 -1711 3222
rect -1745 1214 -1711 1230
rect -1649 3206 -1615 3222
rect -1649 1214 -1615 1230
rect -1553 3206 -1519 3222
rect -1553 1214 -1519 1230
rect -1457 3206 -1423 3222
rect -1457 1214 -1423 1230
rect -1361 3206 -1327 3222
rect -1361 1214 -1327 1230
rect -1265 3206 -1231 3222
rect -1265 1214 -1231 1230
rect -1169 3206 -1135 3222
rect -1169 1214 -1135 1230
rect -1073 3206 -1039 3222
rect -1073 1214 -1039 1230
rect -977 3206 -943 3222
rect -977 1214 -943 1230
rect -881 3206 -847 3222
rect -881 1214 -847 1230
rect -785 3206 -751 3222
rect -785 1214 -751 1230
rect -689 3206 -655 3222
rect -689 1214 -655 1230
rect -593 3206 -559 3222
rect -593 1214 -559 1230
rect -497 3206 -463 3222
rect -497 1214 -463 1230
rect -401 3206 -367 3222
rect -401 1214 -367 1230
rect -305 3206 -271 3222
rect -305 1214 -271 1230
rect -209 3206 -175 3222
rect -209 1214 -175 1230
rect -113 3206 -79 3222
rect -113 1214 -79 1230
rect -17 3206 17 3222
rect -17 1214 17 1230
rect 79 3206 113 3222
rect 79 1214 113 1230
rect 175 3206 209 3222
rect 175 1214 209 1230
rect 271 3206 305 3222
rect 271 1214 305 1230
rect 367 3206 401 3222
rect 367 1214 401 1230
rect 463 3206 497 3222
rect 463 1214 497 1230
rect 559 3206 593 3222
rect 559 1214 593 1230
rect 655 3206 689 3222
rect 655 1214 689 1230
rect 751 3206 785 3222
rect 751 1214 785 1230
rect 847 3206 881 3222
rect 847 1214 881 1230
rect 943 3206 977 3222
rect 943 1214 977 1230
rect 1039 3206 1073 3222
rect 1039 1214 1073 1230
rect 1135 3206 1169 3222
rect 1135 1214 1169 1230
rect 1231 3206 1265 3222
rect 1231 1214 1265 1230
rect 1327 3206 1361 3222
rect 1327 1214 1361 1230
rect 1423 3206 1457 3222
rect 1423 1214 1457 1230
rect 1519 3206 1553 3222
rect 1519 1214 1553 1230
rect 1615 3206 1649 3222
rect 1615 1214 1649 1230
rect 1711 3206 1745 3222
rect 1711 1214 1745 1230
rect 1807 3206 1841 3222
rect 1807 1214 1841 1230
rect 1903 3206 1937 3222
rect 1903 1214 1937 1230
rect 1999 3206 2033 3222
rect 1999 1214 2033 1230
rect 2095 3206 2129 3222
rect 2095 1214 2129 1230
rect 2191 3206 2225 3222
rect 2191 1214 2225 1230
rect 2287 3206 2321 3222
rect 2287 1214 2321 1230
rect 2383 3206 2417 3222
rect 2383 1214 2417 1230
rect 2479 3206 2513 3222
rect 2479 1214 2513 1230
rect 2575 3206 2609 3222
rect 2575 1214 2609 1230
rect 2671 3206 2705 3222
rect 2671 1214 2705 1230
rect 2767 3206 2801 3222
rect 2767 1214 2801 1230
rect 2863 3206 2897 3222
rect 2863 1214 2897 1230
rect -2865 1146 -2849 1180
rect -2815 1146 -2799 1180
rect -2673 1146 -2657 1180
rect -2623 1146 -2607 1180
rect -2481 1146 -2465 1180
rect -2431 1146 -2415 1180
rect -2289 1146 -2273 1180
rect -2239 1146 -2223 1180
rect -2097 1146 -2081 1180
rect -2047 1146 -2031 1180
rect -1905 1146 -1889 1180
rect -1855 1146 -1839 1180
rect -1713 1146 -1697 1180
rect -1663 1146 -1647 1180
rect -1521 1146 -1505 1180
rect -1471 1146 -1455 1180
rect -1329 1146 -1313 1180
rect -1279 1146 -1263 1180
rect -1137 1146 -1121 1180
rect -1087 1146 -1071 1180
rect -945 1146 -929 1180
rect -895 1146 -879 1180
rect -753 1146 -737 1180
rect -703 1146 -687 1180
rect -561 1146 -545 1180
rect -511 1146 -495 1180
rect -369 1146 -353 1180
rect -319 1146 -303 1180
rect -177 1146 -161 1180
rect -127 1146 -111 1180
rect 15 1146 31 1180
rect 65 1146 81 1180
rect 207 1146 223 1180
rect 257 1146 273 1180
rect 399 1146 415 1180
rect 449 1146 465 1180
rect 591 1146 607 1180
rect 641 1146 657 1180
rect 783 1146 799 1180
rect 833 1146 849 1180
rect 975 1146 991 1180
rect 1025 1146 1041 1180
rect 1167 1146 1183 1180
rect 1217 1146 1233 1180
rect 1359 1146 1375 1180
rect 1409 1146 1425 1180
rect 1551 1146 1567 1180
rect 1601 1146 1617 1180
rect 1743 1146 1759 1180
rect 1793 1146 1809 1180
rect 1935 1146 1951 1180
rect 1985 1146 2001 1180
rect 2127 1146 2143 1180
rect 2177 1146 2193 1180
rect 2319 1146 2335 1180
rect 2369 1146 2385 1180
rect 2511 1146 2527 1180
rect 2561 1146 2577 1180
rect 2703 1146 2719 1180
rect 2753 1146 2769 1180
rect -2865 1038 -2849 1072
rect -2815 1038 -2799 1072
rect -2673 1038 -2657 1072
rect -2623 1038 -2607 1072
rect -2481 1038 -2465 1072
rect -2431 1038 -2415 1072
rect -2289 1038 -2273 1072
rect -2239 1038 -2223 1072
rect -2097 1038 -2081 1072
rect -2047 1038 -2031 1072
rect -1905 1038 -1889 1072
rect -1855 1038 -1839 1072
rect -1713 1038 -1697 1072
rect -1663 1038 -1647 1072
rect -1521 1038 -1505 1072
rect -1471 1038 -1455 1072
rect -1329 1038 -1313 1072
rect -1279 1038 -1263 1072
rect -1137 1038 -1121 1072
rect -1087 1038 -1071 1072
rect -945 1038 -929 1072
rect -895 1038 -879 1072
rect -753 1038 -737 1072
rect -703 1038 -687 1072
rect -561 1038 -545 1072
rect -511 1038 -495 1072
rect -369 1038 -353 1072
rect -319 1038 -303 1072
rect -177 1038 -161 1072
rect -127 1038 -111 1072
rect 15 1038 31 1072
rect 65 1038 81 1072
rect 207 1038 223 1072
rect 257 1038 273 1072
rect 399 1038 415 1072
rect 449 1038 465 1072
rect 591 1038 607 1072
rect 641 1038 657 1072
rect 783 1038 799 1072
rect 833 1038 849 1072
rect 975 1038 991 1072
rect 1025 1038 1041 1072
rect 1167 1038 1183 1072
rect 1217 1038 1233 1072
rect 1359 1038 1375 1072
rect 1409 1038 1425 1072
rect 1551 1038 1567 1072
rect 1601 1038 1617 1072
rect 1743 1038 1759 1072
rect 1793 1038 1809 1072
rect 1935 1038 1951 1072
rect 1985 1038 2001 1072
rect 2127 1038 2143 1072
rect 2177 1038 2193 1072
rect 2319 1038 2335 1072
rect 2369 1038 2385 1072
rect 2511 1038 2527 1072
rect 2561 1038 2577 1072
rect 2703 1038 2719 1072
rect 2753 1038 2769 1072
rect -2897 988 -2863 1004
rect -2897 -1004 -2863 -988
rect -2801 988 -2767 1004
rect -2801 -1004 -2767 -988
rect -2705 988 -2671 1004
rect -2705 -1004 -2671 -988
rect -2609 988 -2575 1004
rect -2609 -1004 -2575 -988
rect -2513 988 -2479 1004
rect -2513 -1004 -2479 -988
rect -2417 988 -2383 1004
rect -2417 -1004 -2383 -988
rect -2321 988 -2287 1004
rect -2321 -1004 -2287 -988
rect -2225 988 -2191 1004
rect -2225 -1004 -2191 -988
rect -2129 988 -2095 1004
rect -2129 -1004 -2095 -988
rect -2033 988 -1999 1004
rect -2033 -1004 -1999 -988
rect -1937 988 -1903 1004
rect -1937 -1004 -1903 -988
rect -1841 988 -1807 1004
rect -1841 -1004 -1807 -988
rect -1745 988 -1711 1004
rect -1745 -1004 -1711 -988
rect -1649 988 -1615 1004
rect -1649 -1004 -1615 -988
rect -1553 988 -1519 1004
rect -1553 -1004 -1519 -988
rect -1457 988 -1423 1004
rect -1457 -1004 -1423 -988
rect -1361 988 -1327 1004
rect -1361 -1004 -1327 -988
rect -1265 988 -1231 1004
rect -1265 -1004 -1231 -988
rect -1169 988 -1135 1004
rect -1169 -1004 -1135 -988
rect -1073 988 -1039 1004
rect -1073 -1004 -1039 -988
rect -977 988 -943 1004
rect -977 -1004 -943 -988
rect -881 988 -847 1004
rect -881 -1004 -847 -988
rect -785 988 -751 1004
rect -785 -1004 -751 -988
rect -689 988 -655 1004
rect -689 -1004 -655 -988
rect -593 988 -559 1004
rect -593 -1004 -559 -988
rect -497 988 -463 1004
rect -497 -1004 -463 -988
rect -401 988 -367 1004
rect -401 -1004 -367 -988
rect -305 988 -271 1004
rect -305 -1004 -271 -988
rect -209 988 -175 1004
rect -209 -1004 -175 -988
rect -113 988 -79 1004
rect -113 -1004 -79 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 79 988 113 1004
rect 79 -1004 113 -988
rect 175 988 209 1004
rect 175 -1004 209 -988
rect 271 988 305 1004
rect 271 -1004 305 -988
rect 367 988 401 1004
rect 367 -1004 401 -988
rect 463 988 497 1004
rect 463 -1004 497 -988
rect 559 988 593 1004
rect 559 -1004 593 -988
rect 655 988 689 1004
rect 655 -1004 689 -988
rect 751 988 785 1004
rect 751 -1004 785 -988
rect 847 988 881 1004
rect 847 -1004 881 -988
rect 943 988 977 1004
rect 943 -1004 977 -988
rect 1039 988 1073 1004
rect 1039 -1004 1073 -988
rect 1135 988 1169 1004
rect 1135 -1004 1169 -988
rect 1231 988 1265 1004
rect 1231 -1004 1265 -988
rect 1327 988 1361 1004
rect 1327 -1004 1361 -988
rect 1423 988 1457 1004
rect 1423 -1004 1457 -988
rect 1519 988 1553 1004
rect 1519 -1004 1553 -988
rect 1615 988 1649 1004
rect 1615 -1004 1649 -988
rect 1711 988 1745 1004
rect 1711 -1004 1745 -988
rect 1807 988 1841 1004
rect 1807 -1004 1841 -988
rect 1903 988 1937 1004
rect 1903 -1004 1937 -988
rect 1999 988 2033 1004
rect 1999 -1004 2033 -988
rect 2095 988 2129 1004
rect 2095 -1004 2129 -988
rect 2191 988 2225 1004
rect 2191 -1004 2225 -988
rect 2287 988 2321 1004
rect 2287 -1004 2321 -988
rect 2383 988 2417 1004
rect 2383 -1004 2417 -988
rect 2479 988 2513 1004
rect 2479 -1004 2513 -988
rect 2575 988 2609 1004
rect 2575 -1004 2609 -988
rect 2671 988 2705 1004
rect 2671 -1004 2705 -988
rect 2767 988 2801 1004
rect 2767 -1004 2801 -988
rect 2863 988 2897 1004
rect 2863 -1004 2897 -988
rect -2769 -1072 -2753 -1038
rect -2719 -1072 -2703 -1038
rect -2577 -1072 -2561 -1038
rect -2527 -1072 -2511 -1038
rect -2385 -1072 -2369 -1038
rect -2335 -1072 -2319 -1038
rect -2193 -1072 -2177 -1038
rect -2143 -1072 -2127 -1038
rect -2001 -1072 -1985 -1038
rect -1951 -1072 -1935 -1038
rect -1809 -1072 -1793 -1038
rect -1759 -1072 -1743 -1038
rect -1617 -1072 -1601 -1038
rect -1567 -1072 -1551 -1038
rect -1425 -1072 -1409 -1038
rect -1375 -1072 -1359 -1038
rect -1233 -1072 -1217 -1038
rect -1183 -1072 -1167 -1038
rect -1041 -1072 -1025 -1038
rect -991 -1072 -975 -1038
rect -849 -1072 -833 -1038
rect -799 -1072 -783 -1038
rect -657 -1072 -641 -1038
rect -607 -1072 -591 -1038
rect -465 -1072 -449 -1038
rect -415 -1072 -399 -1038
rect -273 -1072 -257 -1038
rect -223 -1072 -207 -1038
rect -81 -1072 -65 -1038
rect -31 -1072 -15 -1038
rect 111 -1072 127 -1038
rect 161 -1072 177 -1038
rect 303 -1072 319 -1038
rect 353 -1072 369 -1038
rect 495 -1072 511 -1038
rect 545 -1072 561 -1038
rect 687 -1072 703 -1038
rect 737 -1072 753 -1038
rect 879 -1072 895 -1038
rect 929 -1072 945 -1038
rect 1071 -1072 1087 -1038
rect 1121 -1072 1137 -1038
rect 1263 -1072 1279 -1038
rect 1313 -1072 1329 -1038
rect 1455 -1072 1471 -1038
rect 1505 -1072 1521 -1038
rect 1647 -1072 1663 -1038
rect 1697 -1072 1713 -1038
rect 1839 -1072 1855 -1038
rect 1889 -1072 1905 -1038
rect 2031 -1072 2047 -1038
rect 2081 -1072 2097 -1038
rect 2223 -1072 2239 -1038
rect 2273 -1072 2289 -1038
rect 2415 -1072 2431 -1038
rect 2465 -1072 2481 -1038
rect 2607 -1072 2623 -1038
rect 2657 -1072 2673 -1038
rect 2799 -1072 2815 -1038
rect 2849 -1072 2865 -1038
rect -2769 -1180 -2753 -1146
rect -2719 -1180 -2703 -1146
rect -2577 -1180 -2561 -1146
rect -2527 -1180 -2511 -1146
rect -2385 -1180 -2369 -1146
rect -2335 -1180 -2319 -1146
rect -2193 -1180 -2177 -1146
rect -2143 -1180 -2127 -1146
rect -2001 -1180 -1985 -1146
rect -1951 -1180 -1935 -1146
rect -1809 -1180 -1793 -1146
rect -1759 -1180 -1743 -1146
rect -1617 -1180 -1601 -1146
rect -1567 -1180 -1551 -1146
rect -1425 -1180 -1409 -1146
rect -1375 -1180 -1359 -1146
rect -1233 -1180 -1217 -1146
rect -1183 -1180 -1167 -1146
rect -1041 -1180 -1025 -1146
rect -991 -1180 -975 -1146
rect -849 -1180 -833 -1146
rect -799 -1180 -783 -1146
rect -657 -1180 -641 -1146
rect -607 -1180 -591 -1146
rect -465 -1180 -449 -1146
rect -415 -1180 -399 -1146
rect -273 -1180 -257 -1146
rect -223 -1180 -207 -1146
rect -81 -1180 -65 -1146
rect -31 -1180 -15 -1146
rect 111 -1180 127 -1146
rect 161 -1180 177 -1146
rect 303 -1180 319 -1146
rect 353 -1180 369 -1146
rect 495 -1180 511 -1146
rect 545 -1180 561 -1146
rect 687 -1180 703 -1146
rect 737 -1180 753 -1146
rect 879 -1180 895 -1146
rect 929 -1180 945 -1146
rect 1071 -1180 1087 -1146
rect 1121 -1180 1137 -1146
rect 1263 -1180 1279 -1146
rect 1313 -1180 1329 -1146
rect 1455 -1180 1471 -1146
rect 1505 -1180 1521 -1146
rect 1647 -1180 1663 -1146
rect 1697 -1180 1713 -1146
rect 1839 -1180 1855 -1146
rect 1889 -1180 1905 -1146
rect 2031 -1180 2047 -1146
rect 2081 -1180 2097 -1146
rect 2223 -1180 2239 -1146
rect 2273 -1180 2289 -1146
rect 2415 -1180 2431 -1146
rect 2465 -1180 2481 -1146
rect 2607 -1180 2623 -1146
rect 2657 -1180 2673 -1146
rect 2799 -1180 2815 -1146
rect 2849 -1180 2865 -1146
rect -2897 -1230 -2863 -1214
rect -2897 -3222 -2863 -3206
rect -2801 -1230 -2767 -1214
rect -2801 -3222 -2767 -3206
rect -2705 -1230 -2671 -1214
rect -2705 -3222 -2671 -3206
rect -2609 -1230 -2575 -1214
rect -2609 -3222 -2575 -3206
rect -2513 -1230 -2479 -1214
rect -2513 -3222 -2479 -3206
rect -2417 -1230 -2383 -1214
rect -2417 -3222 -2383 -3206
rect -2321 -1230 -2287 -1214
rect -2321 -3222 -2287 -3206
rect -2225 -1230 -2191 -1214
rect -2225 -3222 -2191 -3206
rect -2129 -1230 -2095 -1214
rect -2129 -3222 -2095 -3206
rect -2033 -1230 -1999 -1214
rect -2033 -3222 -1999 -3206
rect -1937 -1230 -1903 -1214
rect -1937 -3222 -1903 -3206
rect -1841 -1230 -1807 -1214
rect -1841 -3222 -1807 -3206
rect -1745 -1230 -1711 -1214
rect -1745 -3222 -1711 -3206
rect -1649 -1230 -1615 -1214
rect -1649 -3222 -1615 -3206
rect -1553 -1230 -1519 -1214
rect -1553 -3222 -1519 -3206
rect -1457 -1230 -1423 -1214
rect -1457 -3222 -1423 -3206
rect -1361 -1230 -1327 -1214
rect -1361 -3222 -1327 -3206
rect -1265 -1230 -1231 -1214
rect -1265 -3222 -1231 -3206
rect -1169 -1230 -1135 -1214
rect -1169 -3222 -1135 -3206
rect -1073 -1230 -1039 -1214
rect -1073 -3222 -1039 -3206
rect -977 -1230 -943 -1214
rect -977 -3222 -943 -3206
rect -881 -1230 -847 -1214
rect -881 -3222 -847 -3206
rect -785 -1230 -751 -1214
rect -785 -3222 -751 -3206
rect -689 -1230 -655 -1214
rect -689 -3222 -655 -3206
rect -593 -1230 -559 -1214
rect -593 -3222 -559 -3206
rect -497 -1230 -463 -1214
rect -497 -3222 -463 -3206
rect -401 -1230 -367 -1214
rect -401 -3222 -367 -3206
rect -305 -1230 -271 -1214
rect -305 -3222 -271 -3206
rect -209 -1230 -175 -1214
rect -209 -3222 -175 -3206
rect -113 -1230 -79 -1214
rect -113 -3222 -79 -3206
rect -17 -1230 17 -1214
rect -17 -3222 17 -3206
rect 79 -1230 113 -1214
rect 79 -3222 113 -3206
rect 175 -1230 209 -1214
rect 175 -3222 209 -3206
rect 271 -1230 305 -1214
rect 271 -3222 305 -3206
rect 367 -1230 401 -1214
rect 367 -3222 401 -3206
rect 463 -1230 497 -1214
rect 463 -3222 497 -3206
rect 559 -1230 593 -1214
rect 559 -3222 593 -3206
rect 655 -1230 689 -1214
rect 655 -3222 689 -3206
rect 751 -1230 785 -1214
rect 751 -3222 785 -3206
rect 847 -1230 881 -1214
rect 847 -3222 881 -3206
rect 943 -1230 977 -1214
rect 943 -3222 977 -3206
rect 1039 -1230 1073 -1214
rect 1039 -3222 1073 -3206
rect 1135 -1230 1169 -1214
rect 1135 -3222 1169 -3206
rect 1231 -1230 1265 -1214
rect 1231 -3222 1265 -3206
rect 1327 -1230 1361 -1214
rect 1327 -3222 1361 -3206
rect 1423 -1230 1457 -1214
rect 1423 -3222 1457 -3206
rect 1519 -1230 1553 -1214
rect 1519 -3222 1553 -3206
rect 1615 -1230 1649 -1214
rect 1615 -3222 1649 -3206
rect 1711 -1230 1745 -1214
rect 1711 -3222 1745 -3206
rect 1807 -1230 1841 -1214
rect 1807 -3222 1841 -3206
rect 1903 -1230 1937 -1214
rect 1903 -3222 1937 -3206
rect 1999 -1230 2033 -1214
rect 1999 -3222 2033 -3206
rect 2095 -1230 2129 -1214
rect 2095 -3222 2129 -3206
rect 2191 -1230 2225 -1214
rect 2191 -3222 2225 -3206
rect 2287 -1230 2321 -1214
rect 2287 -3222 2321 -3206
rect 2383 -1230 2417 -1214
rect 2383 -3222 2417 -3206
rect 2479 -1230 2513 -1214
rect 2479 -3222 2513 -3206
rect 2575 -1230 2609 -1214
rect 2575 -3222 2609 -3206
rect 2671 -1230 2705 -1214
rect 2671 -3222 2705 -3206
rect 2767 -1230 2801 -1214
rect 2767 -3222 2801 -3206
rect 2863 -1230 2897 -1214
rect 2863 -3222 2897 -3206
rect -2865 -3290 -2849 -3256
rect -2815 -3290 -2799 -3256
rect -2673 -3290 -2657 -3256
rect -2623 -3290 -2607 -3256
rect -2481 -3290 -2465 -3256
rect -2431 -3290 -2415 -3256
rect -2289 -3290 -2273 -3256
rect -2239 -3290 -2223 -3256
rect -2097 -3290 -2081 -3256
rect -2047 -3290 -2031 -3256
rect -1905 -3290 -1889 -3256
rect -1855 -3290 -1839 -3256
rect -1713 -3290 -1697 -3256
rect -1663 -3290 -1647 -3256
rect -1521 -3290 -1505 -3256
rect -1471 -3290 -1455 -3256
rect -1329 -3290 -1313 -3256
rect -1279 -3290 -1263 -3256
rect -1137 -3290 -1121 -3256
rect -1087 -3290 -1071 -3256
rect -945 -3290 -929 -3256
rect -895 -3290 -879 -3256
rect -753 -3290 -737 -3256
rect -703 -3290 -687 -3256
rect -561 -3290 -545 -3256
rect -511 -3290 -495 -3256
rect -369 -3290 -353 -3256
rect -319 -3290 -303 -3256
rect -177 -3290 -161 -3256
rect -127 -3290 -111 -3256
rect 15 -3290 31 -3256
rect 65 -3290 81 -3256
rect 207 -3290 223 -3256
rect 257 -3290 273 -3256
rect 399 -3290 415 -3256
rect 449 -3290 465 -3256
rect 591 -3290 607 -3256
rect 641 -3290 657 -3256
rect 783 -3290 799 -3256
rect 833 -3290 849 -3256
rect 975 -3290 991 -3256
rect 1025 -3290 1041 -3256
rect 1167 -3290 1183 -3256
rect 1217 -3290 1233 -3256
rect 1359 -3290 1375 -3256
rect 1409 -3290 1425 -3256
rect 1551 -3290 1567 -3256
rect 1601 -3290 1617 -3256
rect 1743 -3290 1759 -3256
rect 1793 -3290 1809 -3256
rect 1935 -3290 1951 -3256
rect 1985 -3290 2001 -3256
rect 2127 -3290 2143 -3256
rect 2177 -3290 2193 -3256
rect 2319 -3290 2335 -3256
rect 2369 -3290 2385 -3256
rect 2511 -3290 2527 -3256
rect 2561 -3290 2577 -3256
rect 2703 -3290 2719 -3256
rect 2753 -3290 2769 -3256
<< viali >>
rect -2753 3256 -2719 3290
rect -2561 3256 -2527 3290
rect -2369 3256 -2335 3290
rect -2177 3256 -2143 3290
rect -1985 3256 -1951 3290
rect -1793 3256 -1759 3290
rect -1601 3256 -1567 3290
rect -1409 3256 -1375 3290
rect -1217 3256 -1183 3290
rect -1025 3256 -991 3290
rect -833 3256 -799 3290
rect -641 3256 -607 3290
rect -449 3256 -415 3290
rect -257 3256 -223 3290
rect -65 3256 -31 3290
rect 127 3256 161 3290
rect 319 3256 353 3290
rect 511 3256 545 3290
rect 703 3256 737 3290
rect 895 3256 929 3290
rect 1087 3256 1121 3290
rect 1279 3256 1313 3290
rect 1471 3256 1505 3290
rect 1663 3256 1697 3290
rect 1855 3256 1889 3290
rect 2047 3256 2081 3290
rect 2239 3256 2273 3290
rect 2431 3256 2465 3290
rect 2623 3256 2657 3290
rect 2815 3256 2849 3290
rect -2897 1230 -2863 3206
rect -2801 1230 -2767 3206
rect -2705 1230 -2671 3206
rect -2609 1230 -2575 3206
rect -2513 1230 -2479 3206
rect -2417 1230 -2383 3206
rect -2321 1230 -2287 3206
rect -2225 1230 -2191 3206
rect -2129 1230 -2095 3206
rect -2033 1230 -1999 3206
rect -1937 1230 -1903 3206
rect -1841 1230 -1807 3206
rect -1745 1230 -1711 3206
rect -1649 1230 -1615 3206
rect -1553 1230 -1519 3206
rect -1457 1230 -1423 3206
rect -1361 1230 -1327 3206
rect -1265 1230 -1231 3206
rect -1169 1230 -1135 3206
rect -1073 1230 -1039 3206
rect -977 1230 -943 3206
rect -881 1230 -847 3206
rect -785 1230 -751 3206
rect -689 1230 -655 3206
rect -593 1230 -559 3206
rect -497 1230 -463 3206
rect -401 1230 -367 3206
rect -305 1230 -271 3206
rect -209 1230 -175 3206
rect -113 1230 -79 3206
rect -17 1230 17 3206
rect 79 1230 113 3206
rect 175 1230 209 3206
rect 271 1230 305 3206
rect 367 1230 401 3206
rect 463 1230 497 3206
rect 559 1230 593 3206
rect 655 1230 689 3206
rect 751 1230 785 3206
rect 847 1230 881 3206
rect 943 1230 977 3206
rect 1039 1230 1073 3206
rect 1135 1230 1169 3206
rect 1231 1230 1265 3206
rect 1327 1230 1361 3206
rect 1423 1230 1457 3206
rect 1519 1230 1553 3206
rect 1615 1230 1649 3206
rect 1711 1230 1745 3206
rect 1807 1230 1841 3206
rect 1903 1230 1937 3206
rect 1999 1230 2033 3206
rect 2095 1230 2129 3206
rect 2191 1230 2225 3206
rect 2287 1230 2321 3206
rect 2383 1230 2417 3206
rect 2479 1230 2513 3206
rect 2575 1230 2609 3206
rect 2671 1230 2705 3206
rect 2767 1230 2801 3206
rect 2863 1230 2897 3206
rect -2849 1146 -2815 1180
rect -2657 1146 -2623 1180
rect -2465 1146 -2431 1180
rect -2273 1146 -2239 1180
rect -2081 1146 -2047 1180
rect -1889 1146 -1855 1180
rect -1697 1146 -1663 1180
rect -1505 1146 -1471 1180
rect -1313 1146 -1279 1180
rect -1121 1146 -1087 1180
rect -929 1146 -895 1180
rect -737 1146 -703 1180
rect -545 1146 -511 1180
rect -353 1146 -319 1180
rect -161 1146 -127 1180
rect 31 1146 65 1180
rect 223 1146 257 1180
rect 415 1146 449 1180
rect 607 1146 641 1180
rect 799 1146 833 1180
rect 991 1146 1025 1180
rect 1183 1146 1217 1180
rect 1375 1146 1409 1180
rect 1567 1146 1601 1180
rect 1759 1146 1793 1180
rect 1951 1146 1985 1180
rect 2143 1146 2177 1180
rect 2335 1146 2369 1180
rect 2527 1146 2561 1180
rect 2719 1146 2753 1180
rect -2849 1038 -2815 1072
rect -2657 1038 -2623 1072
rect -2465 1038 -2431 1072
rect -2273 1038 -2239 1072
rect -2081 1038 -2047 1072
rect -1889 1038 -1855 1072
rect -1697 1038 -1663 1072
rect -1505 1038 -1471 1072
rect -1313 1038 -1279 1072
rect -1121 1038 -1087 1072
rect -929 1038 -895 1072
rect -737 1038 -703 1072
rect -545 1038 -511 1072
rect -353 1038 -319 1072
rect -161 1038 -127 1072
rect 31 1038 65 1072
rect 223 1038 257 1072
rect 415 1038 449 1072
rect 607 1038 641 1072
rect 799 1038 833 1072
rect 991 1038 1025 1072
rect 1183 1038 1217 1072
rect 1375 1038 1409 1072
rect 1567 1038 1601 1072
rect 1759 1038 1793 1072
rect 1951 1038 1985 1072
rect 2143 1038 2177 1072
rect 2335 1038 2369 1072
rect 2527 1038 2561 1072
rect 2719 1038 2753 1072
rect -2897 -988 -2863 988
rect -2801 -988 -2767 988
rect -2705 -988 -2671 988
rect -2609 -988 -2575 988
rect -2513 -988 -2479 988
rect -2417 -988 -2383 988
rect -2321 -988 -2287 988
rect -2225 -988 -2191 988
rect -2129 -988 -2095 988
rect -2033 -988 -1999 988
rect -1937 -988 -1903 988
rect -1841 -988 -1807 988
rect -1745 -988 -1711 988
rect -1649 -988 -1615 988
rect -1553 -988 -1519 988
rect -1457 -988 -1423 988
rect -1361 -988 -1327 988
rect -1265 -988 -1231 988
rect -1169 -988 -1135 988
rect -1073 -988 -1039 988
rect -977 -988 -943 988
rect -881 -988 -847 988
rect -785 -988 -751 988
rect -689 -988 -655 988
rect -593 -988 -559 988
rect -497 -988 -463 988
rect -401 -988 -367 988
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect 367 -988 401 988
rect 463 -988 497 988
rect 559 -988 593 988
rect 655 -988 689 988
rect 751 -988 785 988
rect 847 -988 881 988
rect 943 -988 977 988
rect 1039 -988 1073 988
rect 1135 -988 1169 988
rect 1231 -988 1265 988
rect 1327 -988 1361 988
rect 1423 -988 1457 988
rect 1519 -988 1553 988
rect 1615 -988 1649 988
rect 1711 -988 1745 988
rect 1807 -988 1841 988
rect 1903 -988 1937 988
rect 1999 -988 2033 988
rect 2095 -988 2129 988
rect 2191 -988 2225 988
rect 2287 -988 2321 988
rect 2383 -988 2417 988
rect 2479 -988 2513 988
rect 2575 -988 2609 988
rect 2671 -988 2705 988
rect 2767 -988 2801 988
rect 2863 -988 2897 988
rect -2753 -1072 -2719 -1038
rect -2561 -1072 -2527 -1038
rect -2369 -1072 -2335 -1038
rect -2177 -1072 -2143 -1038
rect -1985 -1072 -1951 -1038
rect -1793 -1072 -1759 -1038
rect -1601 -1072 -1567 -1038
rect -1409 -1072 -1375 -1038
rect -1217 -1072 -1183 -1038
rect -1025 -1072 -991 -1038
rect -833 -1072 -799 -1038
rect -641 -1072 -607 -1038
rect -449 -1072 -415 -1038
rect -257 -1072 -223 -1038
rect -65 -1072 -31 -1038
rect 127 -1072 161 -1038
rect 319 -1072 353 -1038
rect 511 -1072 545 -1038
rect 703 -1072 737 -1038
rect 895 -1072 929 -1038
rect 1087 -1072 1121 -1038
rect 1279 -1072 1313 -1038
rect 1471 -1072 1505 -1038
rect 1663 -1072 1697 -1038
rect 1855 -1072 1889 -1038
rect 2047 -1072 2081 -1038
rect 2239 -1072 2273 -1038
rect 2431 -1072 2465 -1038
rect 2623 -1072 2657 -1038
rect 2815 -1072 2849 -1038
rect -2753 -1180 -2719 -1146
rect -2561 -1180 -2527 -1146
rect -2369 -1180 -2335 -1146
rect -2177 -1180 -2143 -1146
rect -1985 -1180 -1951 -1146
rect -1793 -1180 -1759 -1146
rect -1601 -1180 -1567 -1146
rect -1409 -1180 -1375 -1146
rect -1217 -1180 -1183 -1146
rect -1025 -1180 -991 -1146
rect -833 -1180 -799 -1146
rect -641 -1180 -607 -1146
rect -449 -1180 -415 -1146
rect -257 -1180 -223 -1146
rect -65 -1180 -31 -1146
rect 127 -1180 161 -1146
rect 319 -1180 353 -1146
rect 511 -1180 545 -1146
rect 703 -1180 737 -1146
rect 895 -1180 929 -1146
rect 1087 -1180 1121 -1146
rect 1279 -1180 1313 -1146
rect 1471 -1180 1505 -1146
rect 1663 -1180 1697 -1146
rect 1855 -1180 1889 -1146
rect 2047 -1180 2081 -1146
rect 2239 -1180 2273 -1146
rect 2431 -1180 2465 -1146
rect 2623 -1180 2657 -1146
rect 2815 -1180 2849 -1146
rect -2897 -3206 -2863 -1230
rect -2801 -3206 -2767 -1230
rect -2705 -3206 -2671 -1230
rect -2609 -3206 -2575 -1230
rect -2513 -3206 -2479 -1230
rect -2417 -3206 -2383 -1230
rect -2321 -3206 -2287 -1230
rect -2225 -3206 -2191 -1230
rect -2129 -3206 -2095 -1230
rect -2033 -3206 -1999 -1230
rect -1937 -3206 -1903 -1230
rect -1841 -3206 -1807 -1230
rect -1745 -3206 -1711 -1230
rect -1649 -3206 -1615 -1230
rect -1553 -3206 -1519 -1230
rect -1457 -3206 -1423 -1230
rect -1361 -3206 -1327 -1230
rect -1265 -3206 -1231 -1230
rect -1169 -3206 -1135 -1230
rect -1073 -3206 -1039 -1230
rect -977 -3206 -943 -1230
rect -881 -3206 -847 -1230
rect -785 -3206 -751 -1230
rect -689 -3206 -655 -1230
rect -593 -3206 -559 -1230
rect -497 -3206 -463 -1230
rect -401 -3206 -367 -1230
rect -305 -3206 -271 -1230
rect -209 -3206 -175 -1230
rect -113 -3206 -79 -1230
rect -17 -3206 17 -1230
rect 79 -3206 113 -1230
rect 175 -3206 209 -1230
rect 271 -3206 305 -1230
rect 367 -3206 401 -1230
rect 463 -3206 497 -1230
rect 559 -3206 593 -1230
rect 655 -3206 689 -1230
rect 751 -3206 785 -1230
rect 847 -3206 881 -1230
rect 943 -3206 977 -1230
rect 1039 -3206 1073 -1230
rect 1135 -3206 1169 -1230
rect 1231 -3206 1265 -1230
rect 1327 -3206 1361 -1230
rect 1423 -3206 1457 -1230
rect 1519 -3206 1553 -1230
rect 1615 -3206 1649 -1230
rect 1711 -3206 1745 -1230
rect 1807 -3206 1841 -1230
rect 1903 -3206 1937 -1230
rect 1999 -3206 2033 -1230
rect 2095 -3206 2129 -1230
rect 2191 -3206 2225 -1230
rect 2287 -3206 2321 -1230
rect 2383 -3206 2417 -1230
rect 2479 -3206 2513 -1230
rect 2575 -3206 2609 -1230
rect 2671 -3206 2705 -1230
rect 2767 -3206 2801 -1230
rect 2863 -3206 2897 -1230
rect -2849 -3290 -2815 -3256
rect -2657 -3290 -2623 -3256
rect -2465 -3290 -2431 -3256
rect -2273 -3290 -2239 -3256
rect -2081 -3290 -2047 -3256
rect -1889 -3290 -1855 -3256
rect -1697 -3290 -1663 -3256
rect -1505 -3290 -1471 -3256
rect -1313 -3290 -1279 -3256
rect -1121 -3290 -1087 -3256
rect -929 -3290 -895 -3256
rect -737 -3290 -703 -3256
rect -545 -3290 -511 -3256
rect -353 -3290 -319 -3256
rect -161 -3290 -127 -3256
rect 31 -3290 65 -3256
rect 223 -3290 257 -3256
rect 415 -3290 449 -3256
rect 607 -3290 641 -3256
rect 799 -3290 833 -3256
rect 991 -3290 1025 -3256
rect 1183 -3290 1217 -3256
rect 1375 -3290 1409 -3256
rect 1567 -3290 1601 -3256
rect 1759 -3290 1793 -3256
rect 1951 -3290 1985 -3256
rect 2143 -3290 2177 -3256
rect 2335 -3290 2369 -3256
rect 2527 -3290 2561 -3256
rect 2719 -3290 2753 -3256
<< metal1 >>
rect -2765 3290 -2707 3296
rect -2765 3256 -2753 3290
rect -2719 3256 -2707 3290
rect -2765 3250 -2707 3256
rect -2573 3290 -2515 3296
rect -2573 3256 -2561 3290
rect -2527 3256 -2515 3290
rect -2573 3250 -2515 3256
rect -2381 3290 -2323 3296
rect -2381 3256 -2369 3290
rect -2335 3256 -2323 3290
rect -2381 3250 -2323 3256
rect -2189 3290 -2131 3296
rect -2189 3256 -2177 3290
rect -2143 3256 -2131 3290
rect -2189 3250 -2131 3256
rect -1997 3290 -1939 3296
rect -1997 3256 -1985 3290
rect -1951 3256 -1939 3290
rect -1997 3250 -1939 3256
rect -1805 3290 -1747 3296
rect -1805 3256 -1793 3290
rect -1759 3256 -1747 3290
rect -1805 3250 -1747 3256
rect -1613 3290 -1555 3296
rect -1613 3256 -1601 3290
rect -1567 3256 -1555 3290
rect -1613 3250 -1555 3256
rect -1421 3290 -1363 3296
rect -1421 3256 -1409 3290
rect -1375 3256 -1363 3290
rect -1421 3250 -1363 3256
rect -1229 3290 -1171 3296
rect -1229 3256 -1217 3290
rect -1183 3256 -1171 3290
rect -1229 3250 -1171 3256
rect -1037 3290 -979 3296
rect -1037 3256 -1025 3290
rect -991 3256 -979 3290
rect -1037 3250 -979 3256
rect -845 3290 -787 3296
rect -845 3256 -833 3290
rect -799 3256 -787 3290
rect -845 3250 -787 3256
rect -653 3290 -595 3296
rect -653 3256 -641 3290
rect -607 3256 -595 3290
rect -653 3250 -595 3256
rect -461 3290 -403 3296
rect -461 3256 -449 3290
rect -415 3256 -403 3290
rect -461 3250 -403 3256
rect -269 3290 -211 3296
rect -269 3256 -257 3290
rect -223 3256 -211 3290
rect -269 3250 -211 3256
rect -77 3290 -19 3296
rect -77 3256 -65 3290
rect -31 3256 -19 3290
rect -77 3250 -19 3256
rect 115 3290 173 3296
rect 115 3256 127 3290
rect 161 3256 173 3290
rect 115 3250 173 3256
rect 307 3290 365 3296
rect 307 3256 319 3290
rect 353 3256 365 3290
rect 307 3250 365 3256
rect 499 3290 557 3296
rect 499 3256 511 3290
rect 545 3256 557 3290
rect 499 3250 557 3256
rect 691 3290 749 3296
rect 691 3256 703 3290
rect 737 3256 749 3290
rect 691 3250 749 3256
rect 883 3290 941 3296
rect 883 3256 895 3290
rect 929 3256 941 3290
rect 883 3250 941 3256
rect 1075 3290 1133 3296
rect 1075 3256 1087 3290
rect 1121 3256 1133 3290
rect 1075 3250 1133 3256
rect 1267 3290 1325 3296
rect 1267 3256 1279 3290
rect 1313 3256 1325 3290
rect 1267 3250 1325 3256
rect 1459 3290 1517 3296
rect 1459 3256 1471 3290
rect 1505 3256 1517 3290
rect 1459 3250 1517 3256
rect 1651 3290 1709 3296
rect 1651 3256 1663 3290
rect 1697 3256 1709 3290
rect 1651 3250 1709 3256
rect 1843 3290 1901 3296
rect 1843 3256 1855 3290
rect 1889 3256 1901 3290
rect 1843 3250 1901 3256
rect 2035 3290 2093 3296
rect 2035 3256 2047 3290
rect 2081 3256 2093 3290
rect 2035 3250 2093 3256
rect 2227 3290 2285 3296
rect 2227 3256 2239 3290
rect 2273 3256 2285 3290
rect 2227 3250 2285 3256
rect 2419 3290 2477 3296
rect 2419 3256 2431 3290
rect 2465 3256 2477 3290
rect 2419 3250 2477 3256
rect 2611 3290 2669 3296
rect 2611 3256 2623 3290
rect 2657 3256 2669 3290
rect 2611 3250 2669 3256
rect 2803 3290 2861 3296
rect 2803 3256 2815 3290
rect 2849 3256 2861 3290
rect 2803 3250 2861 3256
rect -2903 3206 -2857 3218
rect -2903 1230 -2897 3206
rect -2863 1230 -2857 3206
rect -2903 1218 -2857 1230
rect -2807 3206 -2761 3218
rect -2807 1230 -2801 3206
rect -2767 1230 -2761 3206
rect -2807 1218 -2761 1230
rect -2711 3206 -2665 3218
rect -2711 1230 -2705 3206
rect -2671 1230 -2665 3206
rect -2711 1218 -2665 1230
rect -2615 3206 -2569 3218
rect -2615 1230 -2609 3206
rect -2575 1230 -2569 3206
rect -2615 1218 -2569 1230
rect -2519 3206 -2473 3218
rect -2519 1230 -2513 3206
rect -2479 1230 -2473 3206
rect -2519 1218 -2473 1230
rect -2423 3206 -2377 3218
rect -2423 1230 -2417 3206
rect -2383 1230 -2377 3206
rect -2423 1218 -2377 1230
rect -2327 3206 -2281 3218
rect -2327 1230 -2321 3206
rect -2287 1230 -2281 3206
rect -2327 1218 -2281 1230
rect -2231 3206 -2185 3218
rect -2231 1230 -2225 3206
rect -2191 1230 -2185 3206
rect -2231 1218 -2185 1230
rect -2135 3206 -2089 3218
rect -2135 1230 -2129 3206
rect -2095 1230 -2089 3206
rect -2135 1218 -2089 1230
rect -2039 3206 -1993 3218
rect -2039 1230 -2033 3206
rect -1999 1230 -1993 3206
rect -2039 1218 -1993 1230
rect -1943 3206 -1897 3218
rect -1943 1230 -1937 3206
rect -1903 1230 -1897 3206
rect -1943 1218 -1897 1230
rect -1847 3206 -1801 3218
rect -1847 1230 -1841 3206
rect -1807 1230 -1801 3206
rect -1847 1218 -1801 1230
rect -1751 3206 -1705 3218
rect -1751 1230 -1745 3206
rect -1711 1230 -1705 3206
rect -1751 1218 -1705 1230
rect -1655 3206 -1609 3218
rect -1655 1230 -1649 3206
rect -1615 1230 -1609 3206
rect -1655 1218 -1609 1230
rect -1559 3206 -1513 3218
rect -1559 1230 -1553 3206
rect -1519 1230 -1513 3206
rect -1559 1218 -1513 1230
rect -1463 3206 -1417 3218
rect -1463 1230 -1457 3206
rect -1423 1230 -1417 3206
rect -1463 1218 -1417 1230
rect -1367 3206 -1321 3218
rect -1367 1230 -1361 3206
rect -1327 1230 -1321 3206
rect -1367 1218 -1321 1230
rect -1271 3206 -1225 3218
rect -1271 1230 -1265 3206
rect -1231 1230 -1225 3206
rect -1271 1218 -1225 1230
rect -1175 3206 -1129 3218
rect -1175 1230 -1169 3206
rect -1135 1230 -1129 3206
rect -1175 1218 -1129 1230
rect -1079 3206 -1033 3218
rect -1079 1230 -1073 3206
rect -1039 1230 -1033 3206
rect -1079 1218 -1033 1230
rect -983 3206 -937 3218
rect -983 1230 -977 3206
rect -943 1230 -937 3206
rect -983 1218 -937 1230
rect -887 3206 -841 3218
rect -887 1230 -881 3206
rect -847 1230 -841 3206
rect -887 1218 -841 1230
rect -791 3206 -745 3218
rect -791 1230 -785 3206
rect -751 1230 -745 3206
rect -791 1218 -745 1230
rect -695 3206 -649 3218
rect -695 1230 -689 3206
rect -655 1230 -649 3206
rect -695 1218 -649 1230
rect -599 3206 -553 3218
rect -599 1230 -593 3206
rect -559 1230 -553 3206
rect -599 1218 -553 1230
rect -503 3206 -457 3218
rect -503 1230 -497 3206
rect -463 1230 -457 3206
rect -503 1218 -457 1230
rect -407 3206 -361 3218
rect -407 1230 -401 3206
rect -367 1230 -361 3206
rect -407 1218 -361 1230
rect -311 3206 -265 3218
rect -311 1230 -305 3206
rect -271 1230 -265 3206
rect -311 1218 -265 1230
rect -215 3206 -169 3218
rect -215 1230 -209 3206
rect -175 1230 -169 3206
rect -215 1218 -169 1230
rect -119 3206 -73 3218
rect -119 1230 -113 3206
rect -79 1230 -73 3206
rect -119 1218 -73 1230
rect -23 3206 23 3218
rect -23 1230 -17 3206
rect 17 1230 23 3206
rect -23 1218 23 1230
rect 73 3206 119 3218
rect 73 1230 79 3206
rect 113 1230 119 3206
rect 73 1218 119 1230
rect 169 3206 215 3218
rect 169 1230 175 3206
rect 209 1230 215 3206
rect 169 1218 215 1230
rect 265 3206 311 3218
rect 265 1230 271 3206
rect 305 1230 311 3206
rect 265 1218 311 1230
rect 361 3206 407 3218
rect 361 1230 367 3206
rect 401 1230 407 3206
rect 361 1218 407 1230
rect 457 3206 503 3218
rect 457 1230 463 3206
rect 497 1230 503 3206
rect 457 1218 503 1230
rect 553 3206 599 3218
rect 553 1230 559 3206
rect 593 1230 599 3206
rect 553 1218 599 1230
rect 649 3206 695 3218
rect 649 1230 655 3206
rect 689 1230 695 3206
rect 649 1218 695 1230
rect 745 3206 791 3218
rect 745 1230 751 3206
rect 785 1230 791 3206
rect 745 1218 791 1230
rect 841 3206 887 3218
rect 841 1230 847 3206
rect 881 1230 887 3206
rect 841 1218 887 1230
rect 937 3206 983 3218
rect 937 1230 943 3206
rect 977 1230 983 3206
rect 937 1218 983 1230
rect 1033 3206 1079 3218
rect 1033 1230 1039 3206
rect 1073 1230 1079 3206
rect 1033 1218 1079 1230
rect 1129 3206 1175 3218
rect 1129 1230 1135 3206
rect 1169 1230 1175 3206
rect 1129 1218 1175 1230
rect 1225 3206 1271 3218
rect 1225 1230 1231 3206
rect 1265 1230 1271 3206
rect 1225 1218 1271 1230
rect 1321 3206 1367 3218
rect 1321 1230 1327 3206
rect 1361 1230 1367 3206
rect 1321 1218 1367 1230
rect 1417 3206 1463 3218
rect 1417 1230 1423 3206
rect 1457 1230 1463 3206
rect 1417 1218 1463 1230
rect 1513 3206 1559 3218
rect 1513 1230 1519 3206
rect 1553 1230 1559 3206
rect 1513 1218 1559 1230
rect 1609 3206 1655 3218
rect 1609 1230 1615 3206
rect 1649 1230 1655 3206
rect 1609 1218 1655 1230
rect 1705 3206 1751 3218
rect 1705 1230 1711 3206
rect 1745 1230 1751 3206
rect 1705 1218 1751 1230
rect 1801 3206 1847 3218
rect 1801 1230 1807 3206
rect 1841 1230 1847 3206
rect 1801 1218 1847 1230
rect 1897 3206 1943 3218
rect 1897 1230 1903 3206
rect 1937 1230 1943 3206
rect 1897 1218 1943 1230
rect 1993 3206 2039 3218
rect 1993 1230 1999 3206
rect 2033 1230 2039 3206
rect 1993 1218 2039 1230
rect 2089 3206 2135 3218
rect 2089 1230 2095 3206
rect 2129 1230 2135 3206
rect 2089 1218 2135 1230
rect 2185 3206 2231 3218
rect 2185 1230 2191 3206
rect 2225 1230 2231 3206
rect 2185 1218 2231 1230
rect 2281 3206 2327 3218
rect 2281 1230 2287 3206
rect 2321 1230 2327 3206
rect 2281 1218 2327 1230
rect 2377 3206 2423 3218
rect 2377 1230 2383 3206
rect 2417 1230 2423 3206
rect 2377 1218 2423 1230
rect 2473 3206 2519 3218
rect 2473 1230 2479 3206
rect 2513 1230 2519 3206
rect 2473 1218 2519 1230
rect 2569 3206 2615 3218
rect 2569 1230 2575 3206
rect 2609 1230 2615 3206
rect 2569 1218 2615 1230
rect 2665 3206 2711 3218
rect 2665 1230 2671 3206
rect 2705 1230 2711 3206
rect 2665 1218 2711 1230
rect 2761 3206 2807 3218
rect 2761 1230 2767 3206
rect 2801 1230 2807 3206
rect 2761 1218 2807 1230
rect 2857 3206 2903 3218
rect 2857 1230 2863 3206
rect 2897 1230 2903 3206
rect 2857 1218 2903 1230
rect -2861 1180 -2803 1186
rect -2861 1146 -2849 1180
rect -2815 1146 -2803 1180
rect -2861 1140 -2803 1146
rect -2669 1180 -2611 1186
rect -2669 1146 -2657 1180
rect -2623 1146 -2611 1180
rect -2669 1140 -2611 1146
rect -2477 1180 -2419 1186
rect -2477 1146 -2465 1180
rect -2431 1146 -2419 1180
rect -2477 1140 -2419 1146
rect -2285 1180 -2227 1186
rect -2285 1146 -2273 1180
rect -2239 1146 -2227 1180
rect -2285 1140 -2227 1146
rect -2093 1180 -2035 1186
rect -2093 1146 -2081 1180
rect -2047 1146 -2035 1180
rect -2093 1140 -2035 1146
rect -1901 1180 -1843 1186
rect -1901 1146 -1889 1180
rect -1855 1146 -1843 1180
rect -1901 1140 -1843 1146
rect -1709 1180 -1651 1186
rect -1709 1146 -1697 1180
rect -1663 1146 -1651 1180
rect -1709 1140 -1651 1146
rect -1517 1180 -1459 1186
rect -1517 1146 -1505 1180
rect -1471 1146 -1459 1180
rect -1517 1140 -1459 1146
rect -1325 1180 -1267 1186
rect -1325 1146 -1313 1180
rect -1279 1146 -1267 1180
rect -1325 1140 -1267 1146
rect -1133 1180 -1075 1186
rect -1133 1146 -1121 1180
rect -1087 1146 -1075 1180
rect -1133 1140 -1075 1146
rect -941 1180 -883 1186
rect -941 1146 -929 1180
rect -895 1146 -883 1180
rect -941 1140 -883 1146
rect -749 1180 -691 1186
rect -749 1146 -737 1180
rect -703 1146 -691 1180
rect -749 1140 -691 1146
rect -557 1180 -499 1186
rect -557 1146 -545 1180
rect -511 1146 -499 1180
rect -557 1140 -499 1146
rect -365 1180 -307 1186
rect -365 1146 -353 1180
rect -319 1146 -307 1180
rect -365 1140 -307 1146
rect -173 1180 -115 1186
rect -173 1146 -161 1180
rect -127 1146 -115 1180
rect -173 1140 -115 1146
rect 19 1180 77 1186
rect 19 1146 31 1180
rect 65 1146 77 1180
rect 19 1140 77 1146
rect 211 1180 269 1186
rect 211 1146 223 1180
rect 257 1146 269 1180
rect 211 1140 269 1146
rect 403 1180 461 1186
rect 403 1146 415 1180
rect 449 1146 461 1180
rect 403 1140 461 1146
rect 595 1180 653 1186
rect 595 1146 607 1180
rect 641 1146 653 1180
rect 595 1140 653 1146
rect 787 1180 845 1186
rect 787 1146 799 1180
rect 833 1146 845 1180
rect 787 1140 845 1146
rect 979 1180 1037 1186
rect 979 1146 991 1180
rect 1025 1146 1037 1180
rect 979 1140 1037 1146
rect 1171 1180 1229 1186
rect 1171 1146 1183 1180
rect 1217 1146 1229 1180
rect 1171 1140 1229 1146
rect 1363 1180 1421 1186
rect 1363 1146 1375 1180
rect 1409 1146 1421 1180
rect 1363 1140 1421 1146
rect 1555 1180 1613 1186
rect 1555 1146 1567 1180
rect 1601 1146 1613 1180
rect 1555 1140 1613 1146
rect 1747 1180 1805 1186
rect 1747 1146 1759 1180
rect 1793 1146 1805 1180
rect 1747 1140 1805 1146
rect 1939 1180 1997 1186
rect 1939 1146 1951 1180
rect 1985 1146 1997 1180
rect 1939 1140 1997 1146
rect 2131 1180 2189 1186
rect 2131 1146 2143 1180
rect 2177 1146 2189 1180
rect 2131 1140 2189 1146
rect 2323 1180 2381 1186
rect 2323 1146 2335 1180
rect 2369 1146 2381 1180
rect 2323 1140 2381 1146
rect 2515 1180 2573 1186
rect 2515 1146 2527 1180
rect 2561 1146 2573 1180
rect 2515 1140 2573 1146
rect 2707 1180 2765 1186
rect 2707 1146 2719 1180
rect 2753 1146 2765 1180
rect 2707 1140 2765 1146
rect -2861 1072 -2803 1078
rect -2861 1038 -2849 1072
rect -2815 1038 -2803 1072
rect -2861 1032 -2803 1038
rect -2669 1072 -2611 1078
rect -2669 1038 -2657 1072
rect -2623 1038 -2611 1072
rect -2669 1032 -2611 1038
rect -2477 1072 -2419 1078
rect -2477 1038 -2465 1072
rect -2431 1038 -2419 1072
rect -2477 1032 -2419 1038
rect -2285 1072 -2227 1078
rect -2285 1038 -2273 1072
rect -2239 1038 -2227 1072
rect -2285 1032 -2227 1038
rect -2093 1072 -2035 1078
rect -2093 1038 -2081 1072
rect -2047 1038 -2035 1072
rect -2093 1032 -2035 1038
rect -1901 1072 -1843 1078
rect -1901 1038 -1889 1072
rect -1855 1038 -1843 1072
rect -1901 1032 -1843 1038
rect -1709 1072 -1651 1078
rect -1709 1038 -1697 1072
rect -1663 1038 -1651 1072
rect -1709 1032 -1651 1038
rect -1517 1072 -1459 1078
rect -1517 1038 -1505 1072
rect -1471 1038 -1459 1072
rect -1517 1032 -1459 1038
rect -1325 1072 -1267 1078
rect -1325 1038 -1313 1072
rect -1279 1038 -1267 1072
rect -1325 1032 -1267 1038
rect -1133 1072 -1075 1078
rect -1133 1038 -1121 1072
rect -1087 1038 -1075 1072
rect -1133 1032 -1075 1038
rect -941 1072 -883 1078
rect -941 1038 -929 1072
rect -895 1038 -883 1072
rect -941 1032 -883 1038
rect -749 1072 -691 1078
rect -749 1038 -737 1072
rect -703 1038 -691 1072
rect -749 1032 -691 1038
rect -557 1072 -499 1078
rect -557 1038 -545 1072
rect -511 1038 -499 1072
rect -557 1032 -499 1038
rect -365 1072 -307 1078
rect -365 1038 -353 1072
rect -319 1038 -307 1072
rect -365 1032 -307 1038
rect -173 1072 -115 1078
rect -173 1038 -161 1072
rect -127 1038 -115 1072
rect -173 1032 -115 1038
rect 19 1072 77 1078
rect 19 1038 31 1072
rect 65 1038 77 1072
rect 19 1032 77 1038
rect 211 1072 269 1078
rect 211 1038 223 1072
rect 257 1038 269 1072
rect 211 1032 269 1038
rect 403 1072 461 1078
rect 403 1038 415 1072
rect 449 1038 461 1072
rect 403 1032 461 1038
rect 595 1072 653 1078
rect 595 1038 607 1072
rect 641 1038 653 1072
rect 595 1032 653 1038
rect 787 1072 845 1078
rect 787 1038 799 1072
rect 833 1038 845 1072
rect 787 1032 845 1038
rect 979 1072 1037 1078
rect 979 1038 991 1072
rect 1025 1038 1037 1072
rect 979 1032 1037 1038
rect 1171 1072 1229 1078
rect 1171 1038 1183 1072
rect 1217 1038 1229 1072
rect 1171 1032 1229 1038
rect 1363 1072 1421 1078
rect 1363 1038 1375 1072
rect 1409 1038 1421 1072
rect 1363 1032 1421 1038
rect 1555 1072 1613 1078
rect 1555 1038 1567 1072
rect 1601 1038 1613 1072
rect 1555 1032 1613 1038
rect 1747 1072 1805 1078
rect 1747 1038 1759 1072
rect 1793 1038 1805 1072
rect 1747 1032 1805 1038
rect 1939 1072 1997 1078
rect 1939 1038 1951 1072
rect 1985 1038 1997 1072
rect 1939 1032 1997 1038
rect 2131 1072 2189 1078
rect 2131 1038 2143 1072
rect 2177 1038 2189 1072
rect 2131 1032 2189 1038
rect 2323 1072 2381 1078
rect 2323 1038 2335 1072
rect 2369 1038 2381 1072
rect 2323 1032 2381 1038
rect 2515 1072 2573 1078
rect 2515 1038 2527 1072
rect 2561 1038 2573 1072
rect 2515 1032 2573 1038
rect 2707 1072 2765 1078
rect 2707 1038 2719 1072
rect 2753 1038 2765 1072
rect 2707 1032 2765 1038
rect -2903 988 -2857 1000
rect -2903 -988 -2897 988
rect -2863 -988 -2857 988
rect -2903 -1000 -2857 -988
rect -2807 988 -2761 1000
rect -2807 -988 -2801 988
rect -2767 -988 -2761 988
rect -2807 -1000 -2761 -988
rect -2711 988 -2665 1000
rect -2711 -988 -2705 988
rect -2671 -988 -2665 988
rect -2711 -1000 -2665 -988
rect -2615 988 -2569 1000
rect -2615 -988 -2609 988
rect -2575 -988 -2569 988
rect -2615 -1000 -2569 -988
rect -2519 988 -2473 1000
rect -2519 -988 -2513 988
rect -2479 -988 -2473 988
rect -2519 -1000 -2473 -988
rect -2423 988 -2377 1000
rect -2423 -988 -2417 988
rect -2383 -988 -2377 988
rect -2423 -1000 -2377 -988
rect -2327 988 -2281 1000
rect -2327 -988 -2321 988
rect -2287 -988 -2281 988
rect -2327 -1000 -2281 -988
rect -2231 988 -2185 1000
rect -2231 -988 -2225 988
rect -2191 -988 -2185 988
rect -2231 -1000 -2185 -988
rect -2135 988 -2089 1000
rect -2135 -988 -2129 988
rect -2095 -988 -2089 988
rect -2135 -1000 -2089 -988
rect -2039 988 -1993 1000
rect -2039 -988 -2033 988
rect -1999 -988 -1993 988
rect -2039 -1000 -1993 -988
rect -1943 988 -1897 1000
rect -1943 -988 -1937 988
rect -1903 -988 -1897 988
rect -1943 -1000 -1897 -988
rect -1847 988 -1801 1000
rect -1847 -988 -1841 988
rect -1807 -988 -1801 988
rect -1847 -1000 -1801 -988
rect -1751 988 -1705 1000
rect -1751 -988 -1745 988
rect -1711 -988 -1705 988
rect -1751 -1000 -1705 -988
rect -1655 988 -1609 1000
rect -1655 -988 -1649 988
rect -1615 -988 -1609 988
rect -1655 -1000 -1609 -988
rect -1559 988 -1513 1000
rect -1559 -988 -1553 988
rect -1519 -988 -1513 988
rect -1559 -1000 -1513 -988
rect -1463 988 -1417 1000
rect -1463 -988 -1457 988
rect -1423 -988 -1417 988
rect -1463 -1000 -1417 -988
rect -1367 988 -1321 1000
rect -1367 -988 -1361 988
rect -1327 -988 -1321 988
rect -1367 -1000 -1321 -988
rect -1271 988 -1225 1000
rect -1271 -988 -1265 988
rect -1231 -988 -1225 988
rect -1271 -1000 -1225 -988
rect -1175 988 -1129 1000
rect -1175 -988 -1169 988
rect -1135 -988 -1129 988
rect -1175 -1000 -1129 -988
rect -1079 988 -1033 1000
rect -1079 -988 -1073 988
rect -1039 -988 -1033 988
rect -1079 -1000 -1033 -988
rect -983 988 -937 1000
rect -983 -988 -977 988
rect -943 -988 -937 988
rect -983 -1000 -937 -988
rect -887 988 -841 1000
rect -887 -988 -881 988
rect -847 -988 -841 988
rect -887 -1000 -841 -988
rect -791 988 -745 1000
rect -791 -988 -785 988
rect -751 -988 -745 988
rect -791 -1000 -745 -988
rect -695 988 -649 1000
rect -695 -988 -689 988
rect -655 -988 -649 988
rect -695 -1000 -649 -988
rect -599 988 -553 1000
rect -599 -988 -593 988
rect -559 -988 -553 988
rect -599 -1000 -553 -988
rect -503 988 -457 1000
rect -503 -988 -497 988
rect -463 -988 -457 988
rect -503 -1000 -457 -988
rect -407 988 -361 1000
rect -407 -988 -401 988
rect -367 -988 -361 988
rect -407 -1000 -361 -988
rect -311 988 -265 1000
rect -311 -988 -305 988
rect -271 -988 -265 988
rect -311 -1000 -265 -988
rect -215 988 -169 1000
rect -215 -988 -209 988
rect -175 -988 -169 988
rect -215 -1000 -169 -988
rect -119 988 -73 1000
rect -119 -988 -113 988
rect -79 -988 -73 988
rect -119 -1000 -73 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 73 988 119 1000
rect 73 -988 79 988
rect 113 -988 119 988
rect 73 -1000 119 -988
rect 169 988 215 1000
rect 169 -988 175 988
rect 209 -988 215 988
rect 169 -1000 215 -988
rect 265 988 311 1000
rect 265 -988 271 988
rect 305 -988 311 988
rect 265 -1000 311 -988
rect 361 988 407 1000
rect 361 -988 367 988
rect 401 -988 407 988
rect 361 -1000 407 -988
rect 457 988 503 1000
rect 457 -988 463 988
rect 497 -988 503 988
rect 457 -1000 503 -988
rect 553 988 599 1000
rect 553 -988 559 988
rect 593 -988 599 988
rect 553 -1000 599 -988
rect 649 988 695 1000
rect 649 -988 655 988
rect 689 -988 695 988
rect 649 -1000 695 -988
rect 745 988 791 1000
rect 745 -988 751 988
rect 785 -988 791 988
rect 745 -1000 791 -988
rect 841 988 887 1000
rect 841 -988 847 988
rect 881 -988 887 988
rect 841 -1000 887 -988
rect 937 988 983 1000
rect 937 -988 943 988
rect 977 -988 983 988
rect 937 -1000 983 -988
rect 1033 988 1079 1000
rect 1033 -988 1039 988
rect 1073 -988 1079 988
rect 1033 -1000 1079 -988
rect 1129 988 1175 1000
rect 1129 -988 1135 988
rect 1169 -988 1175 988
rect 1129 -1000 1175 -988
rect 1225 988 1271 1000
rect 1225 -988 1231 988
rect 1265 -988 1271 988
rect 1225 -1000 1271 -988
rect 1321 988 1367 1000
rect 1321 -988 1327 988
rect 1361 -988 1367 988
rect 1321 -1000 1367 -988
rect 1417 988 1463 1000
rect 1417 -988 1423 988
rect 1457 -988 1463 988
rect 1417 -1000 1463 -988
rect 1513 988 1559 1000
rect 1513 -988 1519 988
rect 1553 -988 1559 988
rect 1513 -1000 1559 -988
rect 1609 988 1655 1000
rect 1609 -988 1615 988
rect 1649 -988 1655 988
rect 1609 -1000 1655 -988
rect 1705 988 1751 1000
rect 1705 -988 1711 988
rect 1745 -988 1751 988
rect 1705 -1000 1751 -988
rect 1801 988 1847 1000
rect 1801 -988 1807 988
rect 1841 -988 1847 988
rect 1801 -1000 1847 -988
rect 1897 988 1943 1000
rect 1897 -988 1903 988
rect 1937 -988 1943 988
rect 1897 -1000 1943 -988
rect 1993 988 2039 1000
rect 1993 -988 1999 988
rect 2033 -988 2039 988
rect 1993 -1000 2039 -988
rect 2089 988 2135 1000
rect 2089 -988 2095 988
rect 2129 -988 2135 988
rect 2089 -1000 2135 -988
rect 2185 988 2231 1000
rect 2185 -988 2191 988
rect 2225 -988 2231 988
rect 2185 -1000 2231 -988
rect 2281 988 2327 1000
rect 2281 -988 2287 988
rect 2321 -988 2327 988
rect 2281 -1000 2327 -988
rect 2377 988 2423 1000
rect 2377 -988 2383 988
rect 2417 -988 2423 988
rect 2377 -1000 2423 -988
rect 2473 988 2519 1000
rect 2473 -988 2479 988
rect 2513 -988 2519 988
rect 2473 -1000 2519 -988
rect 2569 988 2615 1000
rect 2569 -988 2575 988
rect 2609 -988 2615 988
rect 2569 -1000 2615 -988
rect 2665 988 2711 1000
rect 2665 -988 2671 988
rect 2705 -988 2711 988
rect 2665 -1000 2711 -988
rect 2761 988 2807 1000
rect 2761 -988 2767 988
rect 2801 -988 2807 988
rect 2761 -1000 2807 -988
rect 2857 988 2903 1000
rect 2857 -988 2863 988
rect 2897 -988 2903 988
rect 2857 -1000 2903 -988
rect -2765 -1038 -2707 -1032
rect -2765 -1072 -2753 -1038
rect -2719 -1072 -2707 -1038
rect -2765 -1078 -2707 -1072
rect -2573 -1038 -2515 -1032
rect -2573 -1072 -2561 -1038
rect -2527 -1072 -2515 -1038
rect -2573 -1078 -2515 -1072
rect -2381 -1038 -2323 -1032
rect -2381 -1072 -2369 -1038
rect -2335 -1072 -2323 -1038
rect -2381 -1078 -2323 -1072
rect -2189 -1038 -2131 -1032
rect -2189 -1072 -2177 -1038
rect -2143 -1072 -2131 -1038
rect -2189 -1078 -2131 -1072
rect -1997 -1038 -1939 -1032
rect -1997 -1072 -1985 -1038
rect -1951 -1072 -1939 -1038
rect -1997 -1078 -1939 -1072
rect -1805 -1038 -1747 -1032
rect -1805 -1072 -1793 -1038
rect -1759 -1072 -1747 -1038
rect -1805 -1078 -1747 -1072
rect -1613 -1038 -1555 -1032
rect -1613 -1072 -1601 -1038
rect -1567 -1072 -1555 -1038
rect -1613 -1078 -1555 -1072
rect -1421 -1038 -1363 -1032
rect -1421 -1072 -1409 -1038
rect -1375 -1072 -1363 -1038
rect -1421 -1078 -1363 -1072
rect -1229 -1038 -1171 -1032
rect -1229 -1072 -1217 -1038
rect -1183 -1072 -1171 -1038
rect -1229 -1078 -1171 -1072
rect -1037 -1038 -979 -1032
rect -1037 -1072 -1025 -1038
rect -991 -1072 -979 -1038
rect -1037 -1078 -979 -1072
rect -845 -1038 -787 -1032
rect -845 -1072 -833 -1038
rect -799 -1072 -787 -1038
rect -845 -1078 -787 -1072
rect -653 -1038 -595 -1032
rect -653 -1072 -641 -1038
rect -607 -1072 -595 -1038
rect -653 -1078 -595 -1072
rect -461 -1038 -403 -1032
rect -461 -1072 -449 -1038
rect -415 -1072 -403 -1038
rect -461 -1078 -403 -1072
rect -269 -1038 -211 -1032
rect -269 -1072 -257 -1038
rect -223 -1072 -211 -1038
rect -269 -1078 -211 -1072
rect -77 -1038 -19 -1032
rect -77 -1072 -65 -1038
rect -31 -1072 -19 -1038
rect -77 -1078 -19 -1072
rect 115 -1038 173 -1032
rect 115 -1072 127 -1038
rect 161 -1072 173 -1038
rect 115 -1078 173 -1072
rect 307 -1038 365 -1032
rect 307 -1072 319 -1038
rect 353 -1072 365 -1038
rect 307 -1078 365 -1072
rect 499 -1038 557 -1032
rect 499 -1072 511 -1038
rect 545 -1072 557 -1038
rect 499 -1078 557 -1072
rect 691 -1038 749 -1032
rect 691 -1072 703 -1038
rect 737 -1072 749 -1038
rect 691 -1078 749 -1072
rect 883 -1038 941 -1032
rect 883 -1072 895 -1038
rect 929 -1072 941 -1038
rect 883 -1078 941 -1072
rect 1075 -1038 1133 -1032
rect 1075 -1072 1087 -1038
rect 1121 -1072 1133 -1038
rect 1075 -1078 1133 -1072
rect 1267 -1038 1325 -1032
rect 1267 -1072 1279 -1038
rect 1313 -1072 1325 -1038
rect 1267 -1078 1325 -1072
rect 1459 -1038 1517 -1032
rect 1459 -1072 1471 -1038
rect 1505 -1072 1517 -1038
rect 1459 -1078 1517 -1072
rect 1651 -1038 1709 -1032
rect 1651 -1072 1663 -1038
rect 1697 -1072 1709 -1038
rect 1651 -1078 1709 -1072
rect 1843 -1038 1901 -1032
rect 1843 -1072 1855 -1038
rect 1889 -1072 1901 -1038
rect 1843 -1078 1901 -1072
rect 2035 -1038 2093 -1032
rect 2035 -1072 2047 -1038
rect 2081 -1072 2093 -1038
rect 2035 -1078 2093 -1072
rect 2227 -1038 2285 -1032
rect 2227 -1072 2239 -1038
rect 2273 -1072 2285 -1038
rect 2227 -1078 2285 -1072
rect 2419 -1038 2477 -1032
rect 2419 -1072 2431 -1038
rect 2465 -1072 2477 -1038
rect 2419 -1078 2477 -1072
rect 2611 -1038 2669 -1032
rect 2611 -1072 2623 -1038
rect 2657 -1072 2669 -1038
rect 2611 -1078 2669 -1072
rect 2803 -1038 2861 -1032
rect 2803 -1072 2815 -1038
rect 2849 -1072 2861 -1038
rect 2803 -1078 2861 -1072
rect -2765 -1146 -2707 -1140
rect -2765 -1180 -2753 -1146
rect -2719 -1180 -2707 -1146
rect -2765 -1186 -2707 -1180
rect -2573 -1146 -2515 -1140
rect -2573 -1180 -2561 -1146
rect -2527 -1180 -2515 -1146
rect -2573 -1186 -2515 -1180
rect -2381 -1146 -2323 -1140
rect -2381 -1180 -2369 -1146
rect -2335 -1180 -2323 -1146
rect -2381 -1186 -2323 -1180
rect -2189 -1146 -2131 -1140
rect -2189 -1180 -2177 -1146
rect -2143 -1180 -2131 -1146
rect -2189 -1186 -2131 -1180
rect -1997 -1146 -1939 -1140
rect -1997 -1180 -1985 -1146
rect -1951 -1180 -1939 -1146
rect -1997 -1186 -1939 -1180
rect -1805 -1146 -1747 -1140
rect -1805 -1180 -1793 -1146
rect -1759 -1180 -1747 -1146
rect -1805 -1186 -1747 -1180
rect -1613 -1146 -1555 -1140
rect -1613 -1180 -1601 -1146
rect -1567 -1180 -1555 -1146
rect -1613 -1186 -1555 -1180
rect -1421 -1146 -1363 -1140
rect -1421 -1180 -1409 -1146
rect -1375 -1180 -1363 -1146
rect -1421 -1186 -1363 -1180
rect -1229 -1146 -1171 -1140
rect -1229 -1180 -1217 -1146
rect -1183 -1180 -1171 -1146
rect -1229 -1186 -1171 -1180
rect -1037 -1146 -979 -1140
rect -1037 -1180 -1025 -1146
rect -991 -1180 -979 -1146
rect -1037 -1186 -979 -1180
rect -845 -1146 -787 -1140
rect -845 -1180 -833 -1146
rect -799 -1180 -787 -1146
rect -845 -1186 -787 -1180
rect -653 -1146 -595 -1140
rect -653 -1180 -641 -1146
rect -607 -1180 -595 -1146
rect -653 -1186 -595 -1180
rect -461 -1146 -403 -1140
rect -461 -1180 -449 -1146
rect -415 -1180 -403 -1146
rect -461 -1186 -403 -1180
rect -269 -1146 -211 -1140
rect -269 -1180 -257 -1146
rect -223 -1180 -211 -1146
rect -269 -1186 -211 -1180
rect -77 -1146 -19 -1140
rect -77 -1180 -65 -1146
rect -31 -1180 -19 -1146
rect -77 -1186 -19 -1180
rect 115 -1146 173 -1140
rect 115 -1180 127 -1146
rect 161 -1180 173 -1146
rect 115 -1186 173 -1180
rect 307 -1146 365 -1140
rect 307 -1180 319 -1146
rect 353 -1180 365 -1146
rect 307 -1186 365 -1180
rect 499 -1146 557 -1140
rect 499 -1180 511 -1146
rect 545 -1180 557 -1146
rect 499 -1186 557 -1180
rect 691 -1146 749 -1140
rect 691 -1180 703 -1146
rect 737 -1180 749 -1146
rect 691 -1186 749 -1180
rect 883 -1146 941 -1140
rect 883 -1180 895 -1146
rect 929 -1180 941 -1146
rect 883 -1186 941 -1180
rect 1075 -1146 1133 -1140
rect 1075 -1180 1087 -1146
rect 1121 -1180 1133 -1146
rect 1075 -1186 1133 -1180
rect 1267 -1146 1325 -1140
rect 1267 -1180 1279 -1146
rect 1313 -1180 1325 -1146
rect 1267 -1186 1325 -1180
rect 1459 -1146 1517 -1140
rect 1459 -1180 1471 -1146
rect 1505 -1180 1517 -1146
rect 1459 -1186 1517 -1180
rect 1651 -1146 1709 -1140
rect 1651 -1180 1663 -1146
rect 1697 -1180 1709 -1146
rect 1651 -1186 1709 -1180
rect 1843 -1146 1901 -1140
rect 1843 -1180 1855 -1146
rect 1889 -1180 1901 -1146
rect 1843 -1186 1901 -1180
rect 2035 -1146 2093 -1140
rect 2035 -1180 2047 -1146
rect 2081 -1180 2093 -1146
rect 2035 -1186 2093 -1180
rect 2227 -1146 2285 -1140
rect 2227 -1180 2239 -1146
rect 2273 -1180 2285 -1146
rect 2227 -1186 2285 -1180
rect 2419 -1146 2477 -1140
rect 2419 -1180 2431 -1146
rect 2465 -1180 2477 -1146
rect 2419 -1186 2477 -1180
rect 2611 -1146 2669 -1140
rect 2611 -1180 2623 -1146
rect 2657 -1180 2669 -1146
rect 2611 -1186 2669 -1180
rect 2803 -1146 2861 -1140
rect 2803 -1180 2815 -1146
rect 2849 -1180 2861 -1146
rect 2803 -1186 2861 -1180
rect -2903 -1230 -2857 -1218
rect -2903 -3206 -2897 -1230
rect -2863 -3206 -2857 -1230
rect -2903 -3218 -2857 -3206
rect -2807 -1230 -2761 -1218
rect -2807 -3206 -2801 -1230
rect -2767 -3206 -2761 -1230
rect -2807 -3218 -2761 -3206
rect -2711 -1230 -2665 -1218
rect -2711 -3206 -2705 -1230
rect -2671 -3206 -2665 -1230
rect -2711 -3218 -2665 -3206
rect -2615 -1230 -2569 -1218
rect -2615 -3206 -2609 -1230
rect -2575 -3206 -2569 -1230
rect -2615 -3218 -2569 -3206
rect -2519 -1230 -2473 -1218
rect -2519 -3206 -2513 -1230
rect -2479 -3206 -2473 -1230
rect -2519 -3218 -2473 -3206
rect -2423 -1230 -2377 -1218
rect -2423 -3206 -2417 -1230
rect -2383 -3206 -2377 -1230
rect -2423 -3218 -2377 -3206
rect -2327 -1230 -2281 -1218
rect -2327 -3206 -2321 -1230
rect -2287 -3206 -2281 -1230
rect -2327 -3218 -2281 -3206
rect -2231 -1230 -2185 -1218
rect -2231 -3206 -2225 -1230
rect -2191 -3206 -2185 -1230
rect -2231 -3218 -2185 -3206
rect -2135 -1230 -2089 -1218
rect -2135 -3206 -2129 -1230
rect -2095 -3206 -2089 -1230
rect -2135 -3218 -2089 -3206
rect -2039 -1230 -1993 -1218
rect -2039 -3206 -2033 -1230
rect -1999 -3206 -1993 -1230
rect -2039 -3218 -1993 -3206
rect -1943 -1230 -1897 -1218
rect -1943 -3206 -1937 -1230
rect -1903 -3206 -1897 -1230
rect -1943 -3218 -1897 -3206
rect -1847 -1230 -1801 -1218
rect -1847 -3206 -1841 -1230
rect -1807 -3206 -1801 -1230
rect -1847 -3218 -1801 -3206
rect -1751 -1230 -1705 -1218
rect -1751 -3206 -1745 -1230
rect -1711 -3206 -1705 -1230
rect -1751 -3218 -1705 -3206
rect -1655 -1230 -1609 -1218
rect -1655 -3206 -1649 -1230
rect -1615 -3206 -1609 -1230
rect -1655 -3218 -1609 -3206
rect -1559 -1230 -1513 -1218
rect -1559 -3206 -1553 -1230
rect -1519 -3206 -1513 -1230
rect -1559 -3218 -1513 -3206
rect -1463 -1230 -1417 -1218
rect -1463 -3206 -1457 -1230
rect -1423 -3206 -1417 -1230
rect -1463 -3218 -1417 -3206
rect -1367 -1230 -1321 -1218
rect -1367 -3206 -1361 -1230
rect -1327 -3206 -1321 -1230
rect -1367 -3218 -1321 -3206
rect -1271 -1230 -1225 -1218
rect -1271 -3206 -1265 -1230
rect -1231 -3206 -1225 -1230
rect -1271 -3218 -1225 -3206
rect -1175 -1230 -1129 -1218
rect -1175 -3206 -1169 -1230
rect -1135 -3206 -1129 -1230
rect -1175 -3218 -1129 -3206
rect -1079 -1230 -1033 -1218
rect -1079 -3206 -1073 -1230
rect -1039 -3206 -1033 -1230
rect -1079 -3218 -1033 -3206
rect -983 -1230 -937 -1218
rect -983 -3206 -977 -1230
rect -943 -3206 -937 -1230
rect -983 -3218 -937 -3206
rect -887 -1230 -841 -1218
rect -887 -3206 -881 -1230
rect -847 -3206 -841 -1230
rect -887 -3218 -841 -3206
rect -791 -1230 -745 -1218
rect -791 -3206 -785 -1230
rect -751 -3206 -745 -1230
rect -791 -3218 -745 -3206
rect -695 -1230 -649 -1218
rect -695 -3206 -689 -1230
rect -655 -3206 -649 -1230
rect -695 -3218 -649 -3206
rect -599 -1230 -553 -1218
rect -599 -3206 -593 -1230
rect -559 -3206 -553 -1230
rect -599 -3218 -553 -3206
rect -503 -1230 -457 -1218
rect -503 -3206 -497 -1230
rect -463 -3206 -457 -1230
rect -503 -3218 -457 -3206
rect -407 -1230 -361 -1218
rect -407 -3206 -401 -1230
rect -367 -3206 -361 -1230
rect -407 -3218 -361 -3206
rect -311 -1230 -265 -1218
rect -311 -3206 -305 -1230
rect -271 -3206 -265 -1230
rect -311 -3218 -265 -3206
rect -215 -1230 -169 -1218
rect -215 -3206 -209 -1230
rect -175 -3206 -169 -1230
rect -215 -3218 -169 -3206
rect -119 -1230 -73 -1218
rect -119 -3206 -113 -1230
rect -79 -3206 -73 -1230
rect -119 -3218 -73 -3206
rect -23 -1230 23 -1218
rect -23 -3206 -17 -1230
rect 17 -3206 23 -1230
rect -23 -3218 23 -3206
rect 73 -1230 119 -1218
rect 73 -3206 79 -1230
rect 113 -3206 119 -1230
rect 73 -3218 119 -3206
rect 169 -1230 215 -1218
rect 169 -3206 175 -1230
rect 209 -3206 215 -1230
rect 169 -3218 215 -3206
rect 265 -1230 311 -1218
rect 265 -3206 271 -1230
rect 305 -3206 311 -1230
rect 265 -3218 311 -3206
rect 361 -1230 407 -1218
rect 361 -3206 367 -1230
rect 401 -3206 407 -1230
rect 361 -3218 407 -3206
rect 457 -1230 503 -1218
rect 457 -3206 463 -1230
rect 497 -3206 503 -1230
rect 457 -3218 503 -3206
rect 553 -1230 599 -1218
rect 553 -3206 559 -1230
rect 593 -3206 599 -1230
rect 553 -3218 599 -3206
rect 649 -1230 695 -1218
rect 649 -3206 655 -1230
rect 689 -3206 695 -1230
rect 649 -3218 695 -3206
rect 745 -1230 791 -1218
rect 745 -3206 751 -1230
rect 785 -3206 791 -1230
rect 745 -3218 791 -3206
rect 841 -1230 887 -1218
rect 841 -3206 847 -1230
rect 881 -3206 887 -1230
rect 841 -3218 887 -3206
rect 937 -1230 983 -1218
rect 937 -3206 943 -1230
rect 977 -3206 983 -1230
rect 937 -3218 983 -3206
rect 1033 -1230 1079 -1218
rect 1033 -3206 1039 -1230
rect 1073 -3206 1079 -1230
rect 1033 -3218 1079 -3206
rect 1129 -1230 1175 -1218
rect 1129 -3206 1135 -1230
rect 1169 -3206 1175 -1230
rect 1129 -3218 1175 -3206
rect 1225 -1230 1271 -1218
rect 1225 -3206 1231 -1230
rect 1265 -3206 1271 -1230
rect 1225 -3218 1271 -3206
rect 1321 -1230 1367 -1218
rect 1321 -3206 1327 -1230
rect 1361 -3206 1367 -1230
rect 1321 -3218 1367 -3206
rect 1417 -1230 1463 -1218
rect 1417 -3206 1423 -1230
rect 1457 -3206 1463 -1230
rect 1417 -3218 1463 -3206
rect 1513 -1230 1559 -1218
rect 1513 -3206 1519 -1230
rect 1553 -3206 1559 -1230
rect 1513 -3218 1559 -3206
rect 1609 -1230 1655 -1218
rect 1609 -3206 1615 -1230
rect 1649 -3206 1655 -1230
rect 1609 -3218 1655 -3206
rect 1705 -1230 1751 -1218
rect 1705 -3206 1711 -1230
rect 1745 -3206 1751 -1230
rect 1705 -3218 1751 -3206
rect 1801 -1230 1847 -1218
rect 1801 -3206 1807 -1230
rect 1841 -3206 1847 -1230
rect 1801 -3218 1847 -3206
rect 1897 -1230 1943 -1218
rect 1897 -3206 1903 -1230
rect 1937 -3206 1943 -1230
rect 1897 -3218 1943 -3206
rect 1993 -1230 2039 -1218
rect 1993 -3206 1999 -1230
rect 2033 -3206 2039 -1230
rect 1993 -3218 2039 -3206
rect 2089 -1230 2135 -1218
rect 2089 -3206 2095 -1230
rect 2129 -3206 2135 -1230
rect 2089 -3218 2135 -3206
rect 2185 -1230 2231 -1218
rect 2185 -3206 2191 -1230
rect 2225 -3206 2231 -1230
rect 2185 -3218 2231 -3206
rect 2281 -1230 2327 -1218
rect 2281 -3206 2287 -1230
rect 2321 -3206 2327 -1230
rect 2281 -3218 2327 -3206
rect 2377 -1230 2423 -1218
rect 2377 -3206 2383 -1230
rect 2417 -3206 2423 -1230
rect 2377 -3218 2423 -3206
rect 2473 -1230 2519 -1218
rect 2473 -3206 2479 -1230
rect 2513 -3206 2519 -1230
rect 2473 -3218 2519 -3206
rect 2569 -1230 2615 -1218
rect 2569 -3206 2575 -1230
rect 2609 -3206 2615 -1230
rect 2569 -3218 2615 -3206
rect 2665 -1230 2711 -1218
rect 2665 -3206 2671 -1230
rect 2705 -3206 2711 -1230
rect 2665 -3218 2711 -3206
rect 2761 -1230 2807 -1218
rect 2761 -3206 2767 -1230
rect 2801 -3206 2807 -1230
rect 2761 -3218 2807 -3206
rect 2857 -1230 2903 -1218
rect 2857 -3206 2863 -1230
rect 2897 -3206 2903 -1230
rect 2857 -3218 2903 -3206
rect -2861 -3256 -2803 -3250
rect -2861 -3290 -2849 -3256
rect -2815 -3290 -2803 -3256
rect -2861 -3296 -2803 -3290
rect -2669 -3256 -2611 -3250
rect -2669 -3290 -2657 -3256
rect -2623 -3290 -2611 -3256
rect -2669 -3296 -2611 -3290
rect -2477 -3256 -2419 -3250
rect -2477 -3290 -2465 -3256
rect -2431 -3290 -2419 -3256
rect -2477 -3296 -2419 -3290
rect -2285 -3256 -2227 -3250
rect -2285 -3290 -2273 -3256
rect -2239 -3290 -2227 -3256
rect -2285 -3296 -2227 -3290
rect -2093 -3256 -2035 -3250
rect -2093 -3290 -2081 -3256
rect -2047 -3290 -2035 -3256
rect -2093 -3296 -2035 -3290
rect -1901 -3256 -1843 -3250
rect -1901 -3290 -1889 -3256
rect -1855 -3290 -1843 -3256
rect -1901 -3296 -1843 -3290
rect -1709 -3256 -1651 -3250
rect -1709 -3290 -1697 -3256
rect -1663 -3290 -1651 -3256
rect -1709 -3296 -1651 -3290
rect -1517 -3256 -1459 -3250
rect -1517 -3290 -1505 -3256
rect -1471 -3290 -1459 -3256
rect -1517 -3296 -1459 -3290
rect -1325 -3256 -1267 -3250
rect -1325 -3290 -1313 -3256
rect -1279 -3290 -1267 -3256
rect -1325 -3296 -1267 -3290
rect -1133 -3256 -1075 -3250
rect -1133 -3290 -1121 -3256
rect -1087 -3290 -1075 -3256
rect -1133 -3296 -1075 -3290
rect -941 -3256 -883 -3250
rect -941 -3290 -929 -3256
rect -895 -3290 -883 -3256
rect -941 -3296 -883 -3290
rect -749 -3256 -691 -3250
rect -749 -3290 -737 -3256
rect -703 -3290 -691 -3256
rect -749 -3296 -691 -3290
rect -557 -3256 -499 -3250
rect -557 -3290 -545 -3256
rect -511 -3290 -499 -3256
rect -557 -3296 -499 -3290
rect -365 -3256 -307 -3250
rect -365 -3290 -353 -3256
rect -319 -3290 -307 -3256
rect -365 -3296 -307 -3290
rect -173 -3256 -115 -3250
rect -173 -3290 -161 -3256
rect -127 -3290 -115 -3256
rect -173 -3296 -115 -3290
rect 19 -3256 77 -3250
rect 19 -3290 31 -3256
rect 65 -3290 77 -3256
rect 19 -3296 77 -3290
rect 211 -3256 269 -3250
rect 211 -3290 223 -3256
rect 257 -3290 269 -3256
rect 211 -3296 269 -3290
rect 403 -3256 461 -3250
rect 403 -3290 415 -3256
rect 449 -3290 461 -3256
rect 403 -3296 461 -3290
rect 595 -3256 653 -3250
rect 595 -3290 607 -3256
rect 641 -3290 653 -3256
rect 595 -3296 653 -3290
rect 787 -3256 845 -3250
rect 787 -3290 799 -3256
rect 833 -3290 845 -3256
rect 787 -3296 845 -3290
rect 979 -3256 1037 -3250
rect 979 -3290 991 -3256
rect 1025 -3290 1037 -3256
rect 979 -3296 1037 -3290
rect 1171 -3256 1229 -3250
rect 1171 -3290 1183 -3256
rect 1217 -3290 1229 -3256
rect 1171 -3296 1229 -3290
rect 1363 -3256 1421 -3250
rect 1363 -3290 1375 -3256
rect 1409 -3290 1421 -3256
rect 1363 -3296 1421 -3290
rect 1555 -3256 1613 -3250
rect 1555 -3290 1567 -3256
rect 1601 -3290 1613 -3256
rect 1555 -3296 1613 -3290
rect 1747 -3256 1805 -3250
rect 1747 -3290 1759 -3256
rect 1793 -3290 1805 -3256
rect 1747 -3296 1805 -3290
rect 1939 -3256 1997 -3250
rect 1939 -3290 1951 -3256
rect 1985 -3290 1997 -3256
rect 1939 -3296 1997 -3290
rect 2131 -3256 2189 -3250
rect 2131 -3290 2143 -3256
rect 2177 -3290 2189 -3256
rect 2131 -3296 2189 -3290
rect 2323 -3256 2381 -3250
rect 2323 -3290 2335 -3256
rect 2369 -3290 2381 -3256
rect 2323 -3296 2381 -3290
rect 2515 -3256 2573 -3250
rect 2515 -3290 2527 -3256
rect 2561 -3290 2573 -3256
rect 2515 -3296 2573 -3290
rect 2707 -3256 2765 -3250
rect 2707 -3290 2719 -3256
rect 2753 -3290 2765 -3256
rect 2707 -3296 2765 -3290
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 10 l 0.150 m 3 nf 60 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
