magic
tech sky130A
magscale 1 2
timestamp 1697743316
<< error_s >>
rect 298 1115 333 1149
rect 299 1096 333 1115
rect 129 1047 187 1053
rect 129 1013 141 1047
rect 129 1007 187 1013
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 318 583 333 1096
rect 352 1062 387 1096
rect 667 1062 702 1079
rect 352 583 386 1062
rect 668 1061 702 1062
rect 668 1025 738 1061
rect 498 994 556 1000
rect 498 960 510 994
rect 685 991 756 1025
rect 1036 991 1071 1025
rect 498 954 556 960
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 352 549 367 583
rect 685 530 755 991
rect 1037 972 1071 991
rect 1423 972 1476 973
rect 867 923 925 929
rect 867 889 879 923
rect 867 883 925 889
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 685 494 738 530
rect 1056 477 1071 972
rect 1090 938 1125 972
rect 1405 938 1476 972
rect 1090 477 1124 938
rect 1406 937 1476 938
rect 1423 903 1494 937
rect 1774 903 1809 920
rect 1236 870 1294 876
rect 1236 836 1248 870
rect 1236 830 1294 836
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1090 443 1105 477
rect 1423 424 1493 903
rect 1775 902 1809 903
rect 1775 866 1845 902
rect 1605 835 1663 841
rect 1605 801 1617 835
rect 1792 832 1863 866
rect 1605 795 1663 801
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1423 388 1476 424
rect 1792 371 1862 832
rect 1974 764 2032 770
rect 1974 730 1986 764
rect 1974 724 2032 730
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1792 335 1845 371
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 1695550690
transform 1 0 158 0 1 866
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 1695550690
transform 1 0 527 0 1 813
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM3
timestamp 1695550690
transform 1 0 896 0 1 751
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1695550690
transform 1 0 1265 0 1 698
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM5
timestamp 1695550690
transform 1 0 1634 0 1 654
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM6
timestamp 1695550690
transform 1 0 2003 0 1 592
box -211 -310 211 310
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 A
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 B
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>
