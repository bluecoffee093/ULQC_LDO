magic
tech sky130A
magscale 1 2
timestamp 1695685220
<< error_p >>
rect 560946 696204 561528 696232
<< metal1 >>
rect 70042 588912 71614 696752
rect 70014 587298 227256 588912
rect 229234 588054 230288 699890
rect 249330 671696 249588 671700
rect 318996 671696 323898 697254
rect 560946 696204 561528 696206
rect 560904 677982 579550 682990
rect 249330 671354 323898 671696
rect 249330 593942 249588 671354
rect 318996 669538 323898 671354
rect 560946 646680 561550 677982
rect 251288 646316 561550 646680
rect 251288 646312 561548 646316
rect 249328 593844 249588 593942
rect 249328 588174 249586 593844
rect 250940 592422 250950 592644
rect 251150 592422 251160 592644
rect 70014 587150 224660 587298
rect 224650 587146 224660 587150
rect 227262 587146 227272 587298
rect 229238 586488 230284 588054
rect 249328 587972 250806 588174
rect 247854 587662 250470 587664
rect 247848 587460 247858 587662
rect 248062 587464 250470 587662
rect 250948 587466 251148 592422
rect 251290 592000 251530 646312
rect 253596 613054 253606 616202
rect 253900 613054 253910 616202
rect 253604 612158 253906 613054
rect 251290 591866 251532 592000
rect 251292 587940 251532 591866
rect 252188 590848 252198 591564
rect 252436 590848 252446 591564
rect 252198 587900 252438 590848
rect 248062 587460 248072 587464
rect 250594 587096 250604 587296
rect 250804 587096 250814 587296
rect 251266 587096 251276 587296
rect 251476 587096 251486 587296
rect 253618 587290 253898 612158
rect 570052 593918 570062 594480
rect 570460 593918 570470 594480
rect 258596 593592 259018 593620
rect 258586 593088 258596 593592
rect 259020 593088 259030 593592
rect 251846 587086 251856 587286
rect 252056 587086 252066 587286
rect 252462 587084 252472 587284
rect 252672 587084 252682 587284
rect 252910 587092 253898 587290
rect 253618 587086 253898 587092
rect 248284 586910 250438 586912
rect 248282 586712 250438 586910
rect 229230 586474 247574 586488
rect 229230 586274 247246 586474
rect 247576 586274 247586 586474
rect 229230 586256 247574 586274
rect 79356 585498 79366 585500
rect 51584 585254 79366 585498
rect 79672 585254 79682 585500
rect 51584 564244 57966 585254
rect 17818 559410 57978 564244
rect 51584 559372 57966 559410
rect 61492 536482 61502 536716
rect 61792 536712 61802 536716
rect 61792 536694 72312 536712
rect 61792 536484 71970 536694
rect 72312 536484 72322 536694
rect 61792 536482 61802 536484
rect 10326 499348 10336 500976
rect 12198 500952 12208 500976
rect 75784 500952 75794 500954
rect 12198 499350 75794 500952
rect 78128 499350 78138 500954
rect 12198 499348 12208 499350
rect 248282 474848 248542 586712
rect 249000 586472 250684 586476
rect 248994 586274 249004 586472
rect 249250 586276 250684 586472
rect 249250 586274 249260 586276
rect 250958 585502 251176 586904
rect 253744 586490 253986 586492
rect 253028 586276 255986 586490
rect 250948 585256 250958 585502
rect 251176 585256 251186 585502
rect 248278 311944 248544 474848
rect 248272 311796 248544 311944
rect 248272 168786 248538 311796
rect 253744 197748 253986 586276
rect 258596 585284 259018 593088
rect 570062 590196 570462 593918
rect 570058 589920 570068 590196
rect 570462 589920 570472 590196
rect 570062 589918 570462 589920
rect 258588 585090 258598 585284
rect 259018 585090 259028 585284
rect 258596 585088 259018 585090
rect 253744 197546 567938 197748
rect 253744 197538 253986 197546
rect 565856 181418 567938 197546
rect 572374 168800 574026 168816
rect 572072 168798 574026 168800
rect 519508 168786 574026 168798
rect 248268 168380 574026 168786
rect 519508 168374 574026 168380
rect 572374 136838 574026 168374
<< via1 >>
rect 250950 592422 251150 592644
rect 224660 587146 227262 587298
rect 247858 587460 248062 587662
rect 253606 613054 253900 616202
rect 252198 590848 252436 591564
rect 250604 587096 250804 587296
rect 251276 587096 251476 587296
rect 570062 593918 570460 594480
rect 258596 593088 259020 593592
rect 251856 587086 252056 587286
rect 252472 587084 252672 587284
rect 247246 586274 247576 586474
rect 79366 585254 79672 585500
rect 61502 536482 61792 536716
rect 71970 536484 72312 536694
rect 10336 499348 12198 500976
rect 75794 499350 78128 500954
rect 249004 586274 249250 586472
rect 250958 585256 251176 585502
rect 570068 589920 570462 590196
rect 258598 585090 259018 585284
<< metal2 >>
rect 32758 699214 33394 699280
rect 16202 696096 33394 699214
rect 10390 500986 12190 685176
rect 32758 536716 33394 696096
rect 121900 594118 123554 694480
rect 177234 616562 180314 697868
rect 570062 657162 570456 698566
rect 177118 616208 180320 616562
rect 177118 616202 252734 616208
rect 253606 616202 253900 616212
rect 177118 615898 253606 616202
rect 177140 613076 253606 615898
rect 252470 613064 253606 613076
rect 253900 613064 257426 616202
rect 253606 613044 253900 613054
rect 570064 594490 570456 657162
rect 570062 594480 570460 594490
rect 121814 593602 195218 594118
rect 570062 593908 570460 593918
rect 121814 593592 259020 593602
rect 121814 593088 258596 593592
rect 121814 593086 259020 593088
rect 121814 592296 195218 593086
rect 258596 593078 259020 593086
rect 250950 592644 251150 592654
rect 571898 592644 572242 592646
rect 251150 592422 572242 592644
rect 250950 592412 251150 592422
rect 64902 591564 66344 591576
rect 252198 591564 252436 591574
rect 64902 590848 252198 591564
rect 252436 590848 252450 591564
rect 61502 536716 61792 536726
rect 32236 536484 61502 536716
rect 61502 536472 61792 536482
rect 10336 500976 12198 500986
rect 10336 499338 12198 499348
rect 64902 209704 66344 590848
rect 252198 590838 252436 590848
rect 570068 590200 570462 590206
rect 247854 590196 570462 590200
rect 247854 589926 570068 590196
rect 247858 587662 248062 589926
rect 570068 589910 570462 589920
rect 247858 587450 248062 587460
rect 224660 587298 227262 587308
rect 250604 587296 250804 587306
rect 246604 587294 250604 587296
rect 227262 587146 250604 587294
rect 224660 587136 250604 587146
rect 224662 587098 250604 587136
rect 246604 587096 250604 587098
rect 250604 587086 250804 587096
rect 251276 587296 251476 587306
rect 247246 586474 247576 586484
rect 249004 586474 249250 586482
rect 247576 586472 249250 586474
rect 247576 586274 249004 586472
rect 247246 586264 247576 586274
rect 249004 586264 249250 586274
rect 79366 585502 79672 585510
rect 250958 585502 251176 585512
rect 79366 585500 250958 585502
rect 79672 585256 250958 585500
rect 251276 585488 251476 587096
rect 251856 587286 252056 587296
rect 251856 585534 252056 587086
rect 252472 587284 252672 587294
rect 79366 585244 79672 585254
rect 250958 585246 251176 585256
rect 251280 557614 251474 585488
rect 71970 536694 72312 536704
rect 251280 536694 251476 557614
rect 72312 536484 251476 536694
rect 71970 536478 251476 536484
rect 71970 536474 72312 536478
rect 75794 500960 78128 500964
rect 251854 500960 252058 585534
rect 252472 585280 252672 587084
rect 258598 585284 259018 585294
rect 255232 585280 258598 585282
rect 252460 585098 258598 585280
rect 255232 585094 258598 585098
rect 258598 585080 259018 585090
rect 571898 542534 572242 592422
rect 75782 500954 252198 500960
rect 75782 499350 75794 500954
rect 78128 499350 252198 500954
rect 75782 499312 252198 499350
rect 7640 205064 66344 209704
rect 7640 205032 66294 205064
use ulqc_ldo  ulqc_ldo_0
timestamp 1695554724
transform 1 0 -4393330 0 1 1242836
box 2442 -2542 5374 -645
use user_analog_proj_example  user_analog_proj_example_0 /foss/designs/cass/repo/ULQC_LDO/mag
timestamp 1695673762
transform 1 0 245230 0 1 578608
box 5008 7668 7940 9565
use user_analog_project_wrapper_empty  user_analog_project_wrapper_empty_0 /foss/designs/cass/repo/ULQC_LDO/mag
timestamp 1632839657
transform 1 0 0 0 1 0
box -800 -800 584800 704800
<< end >>
