magic
tech sky130A
magscale 1 2
timestamp 1697926798
<< nmoslvt >>
rect -5261 -3000 -4261 3000
rect -4203 -3000 -3203 3000
rect -3145 -3000 -2145 3000
rect -2087 -3000 -1087 3000
rect -1029 -3000 -29 3000
rect 29 -3000 1029 3000
rect 1087 -3000 2087 3000
rect 2145 -3000 3145 3000
rect 3203 -3000 4203 3000
rect 4261 -3000 5261 3000
<< ndiff >>
rect -5319 2988 -5261 3000
rect -5319 -2988 -5307 2988
rect -5273 -2988 -5261 2988
rect -5319 -3000 -5261 -2988
rect -4261 2988 -4203 3000
rect -4261 -2988 -4249 2988
rect -4215 -2988 -4203 2988
rect -4261 -3000 -4203 -2988
rect -3203 2988 -3145 3000
rect -3203 -2988 -3191 2988
rect -3157 -2988 -3145 2988
rect -3203 -3000 -3145 -2988
rect -2145 2988 -2087 3000
rect -2145 -2988 -2133 2988
rect -2099 -2988 -2087 2988
rect -2145 -3000 -2087 -2988
rect -1087 2988 -1029 3000
rect -1087 -2988 -1075 2988
rect -1041 -2988 -1029 2988
rect -1087 -3000 -1029 -2988
rect -29 2988 29 3000
rect -29 -2988 -17 2988
rect 17 -2988 29 2988
rect -29 -3000 29 -2988
rect 1029 2988 1087 3000
rect 1029 -2988 1041 2988
rect 1075 -2988 1087 2988
rect 1029 -3000 1087 -2988
rect 2087 2988 2145 3000
rect 2087 -2988 2099 2988
rect 2133 -2988 2145 2988
rect 2087 -3000 2145 -2988
rect 3145 2988 3203 3000
rect 3145 -2988 3157 2988
rect 3191 -2988 3203 2988
rect 3145 -3000 3203 -2988
rect 4203 2988 4261 3000
rect 4203 -2988 4215 2988
rect 4249 -2988 4261 2988
rect 4203 -3000 4261 -2988
rect 5261 2988 5319 3000
rect 5261 -2988 5273 2988
rect 5307 -2988 5319 2988
rect 5261 -3000 5319 -2988
<< ndiffc >>
rect -5307 -2988 -5273 2988
rect -4249 -2988 -4215 2988
rect -3191 -2988 -3157 2988
rect -2133 -2988 -2099 2988
rect -1075 -2988 -1041 2988
rect -17 -2988 17 2988
rect 1041 -2988 1075 2988
rect 2099 -2988 2133 2988
rect 3157 -2988 3191 2988
rect 4215 -2988 4249 2988
rect 5273 -2988 5307 2988
<< poly >>
rect -5261 3000 -4261 3026
rect -4203 3000 -3203 3026
rect -3145 3000 -2145 3026
rect -2087 3000 -1087 3026
rect -1029 3000 -29 3026
rect 29 3000 1029 3026
rect 1087 3000 2087 3026
rect 2145 3000 3145 3026
rect 3203 3000 4203 3026
rect 4261 3000 5261 3026
rect -5261 -3026 -4261 -3000
rect -4203 -3026 -3203 -3000
rect -3145 -3026 -2145 -3000
rect -2087 -3026 -1087 -3000
rect -1029 -3026 -29 -3000
rect 29 -3026 1029 -3000
rect 1087 -3026 2087 -3000
rect 2145 -3026 3145 -3000
rect 3203 -3026 4203 -3000
rect 4261 -3026 5261 -3000
<< locali >>
rect -5307 2988 -5273 3004
rect -5307 -3004 -5273 -2988
rect -4249 2988 -4215 3004
rect -4249 -3004 -4215 -2988
rect -3191 2988 -3157 3004
rect -3191 -3004 -3157 -2988
rect -2133 2988 -2099 3004
rect -2133 -3004 -2099 -2988
rect -1075 2988 -1041 3004
rect -1075 -3004 -1041 -2988
rect -17 2988 17 3004
rect -17 -3004 17 -2988
rect 1041 2988 1075 3004
rect 1041 -3004 1075 -2988
rect 2099 2988 2133 3004
rect 2099 -3004 2133 -2988
rect 3157 2988 3191 3004
rect 3157 -3004 3191 -2988
rect 4215 2988 4249 3004
rect 4215 -3004 4249 -2988
rect 5273 2988 5307 3004
rect 5273 -3004 5307 -2988
<< viali >>
rect -5307 -2988 -5273 2988
rect -4249 -2988 -4215 2988
rect -3191 -2988 -3157 2988
rect -2133 -2988 -2099 2988
rect -1075 -2988 -1041 2988
rect -17 -2988 17 2988
rect 1041 -2988 1075 2988
rect 2099 -2988 2133 2988
rect 3157 -2988 3191 2988
rect 4215 -2988 4249 2988
rect 5273 -2988 5307 2988
<< metal1 >>
rect -5313 2988 -5267 3000
rect -5313 -2988 -5307 2988
rect -5273 -2988 -5267 2988
rect -5313 -3000 -5267 -2988
rect -4255 2988 -4209 3000
rect -4255 -2988 -4249 2988
rect -4215 -2988 -4209 2988
rect -4255 -3000 -4209 -2988
rect -3197 2988 -3151 3000
rect -3197 -2988 -3191 2988
rect -3157 -2988 -3151 2988
rect -3197 -3000 -3151 -2988
rect -2139 2988 -2093 3000
rect -2139 -2988 -2133 2988
rect -2099 -2988 -2093 2988
rect -2139 -3000 -2093 -2988
rect -1081 2988 -1035 3000
rect -1081 -2988 -1075 2988
rect -1041 -2988 -1035 2988
rect -1081 -3000 -1035 -2988
rect -23 2988 23 3000
rect -23 -2988 -17 2988
rect 17 -2988 23 2988
rect -23 -3000 23 -2988
rect 1035 2988 1081 3000
rect 1035 -2988 1041 2988
rect 1075 -2988 1081 2988
rect 1035 -3000 1081 -2988
rect 2093 2988 2139 3000
rect 2093 -2988 2099 2988
rect 2133 -2988 2139 2988
rect 2093 -3000 2139 -2988
rect 3151 2988 3197 3000
rect 3151 -2988 3157 2988
rect 3191 -2988 3197 2988
rect 3151 -3000 3197 -2988
rect 4209 2988 4255 3000
rect 4209 -2988 4215 2988
rect 4249 -2988 4255 2988
rect 4209 -3000 4255 -2988
rect 5267 2988 5313 3000
rect 5267 -2988 5273 2988
rect 5307 -2988 5313 2988
rect 5267 -3000 5313 -2988
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 30.0 l 5.0 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
