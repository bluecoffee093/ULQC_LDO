magic
tech sky130A
magscale 1 2
timestamp 1697926267
<< pwell >>
rect -201 -3298 201 3298
<< psubdiff >>
rect -165 3228 -69 3262
rect 69 3228 165 3262
rect -165 3166 -131 3228
rect 131 3166 165 3228
rect -165 -3228 -131 -3166
rect 131 -3228 165 -3166
rect -165 -3262 -69 -3228
rect 69 -3262 165 -3228
<< psubdiffcont >>
rect -69 3228 69 3262
rect -165 -3166 -131 3166
rect 131 -3166 165 3166
rect -69 -3262 69 -3228
<< xpolycontact >>
rect -35 2700 35 3132
rect -35 -3132 35 -2700
<< ppolyres >>
rect -35 -2700 35 2700
<< locali >>
rect -165 3228 -69 3262
rect 69 3228 165 3262
rect -165 3166 -131 3228
rect 131 3166 165 3228
rect -165 -3228 -131 -3166
rect 131 -3228 165 -3166
rect -165 -3262 -69 -3228
rect 69 -3262 165 -3228
<< viali >>
rect -19 2717 19 3114
rect -19 -3114 19 -2717
<< metal1 >>
rect -25 3114 25 3126
rect -25 2717 -19 3114
rect 19 2717 25 3114
rect -25 2705 25 2717
rect -25 -2717 25 -2705
rect -25 -3114 -19 -2717
rect 19 -3114 25 -2717
rect -25 -3126 25 -3114
<< res0p35 >>
rect -37 -2702 37 2702
<< properties >>
string FIXED_BBOX -148 -3245 148 3245
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 27.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 25.783k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
