* SPICE3 file created from user_analog_project_wrapper.ext - technology: sky130A

C0 user_analog_proj_example_0/ulqc_ldo_0/VIN2 user_analog_project_wrapper_empty_0/io_analog[7] 2.05fF
C1 user_analog_project_wrapper_empty_0/io_analog[4] user_analog_project_wrapper_empty_0/io_analog[6] 4.34fF
C2 user_analog_project_wrapper_empty_0/io_analog[0] user_analog_project_wrapper_empty_0/io_analog[1] 10.61fF
C3 user_analog_project_wrapper_empty_0/io_analog[10] user_analog_project_wrapper_empty_0/vssa2 21.81fF
C4 user_analog_project_wrapper_empty_0/io_analog[7] user_analog_project_wrapper_empty_0/vdda2 9.14fF
C5 user_analog_project_wrapper_empty_0/io_analog[5] user_analog_project_wrapper_empty_0/io_analog[6] 13.20fF
C6 user_analog_project_wrapper_empty_0/io_analog[10] user_analog_project_wrapper_empty_0/vdda2 9.85fF
C7 user_analog_project_wrapper_empty_0/io_analog[5] user_analog_project_wrapper_empty_0/vdda2 4.87fF
C8 user_analog_project_wrapper_empty_0/io_analog[10] user_analog_project_wrapper_empty_0/io_analog[9] 4.57fF
C9 user_analog_proj_example_0/ulqc_ldo_0/VIN2 user_analog_project_wrapper_empty_0/io_analog[0] 2.08fF
C10 user_analog_project_wrapper_empty_0/io_analog[8] user_analog_project_wrapper_empty_0/vdda2 6.11fF
C11 user_analog_project_wrapper_empty_0/vssa2 user_analog_project_wrapper_empty_0/vdda2 2.01fF
C12 user_analog_project_wrapper_empty_0/io_analog[0] user_analog_project_wrapper_empty_0/io_analog[6] 4.14fF
C13 user_analog_project_wrapper_empty_0/io_analog[5] user_analog_project_wrapper_empty_0/io_analog[7] 3.06fF
C14 user_analog_project_wrapper_empty_0/vssa2 user_analog_project_wrapper_empty_0/io_analog[9] 14.44fF
C15 user_analog_proj_example_0/ulqc_ldo_0/VIN2 user_analog_project_wrapper_empty_0/io_analog[1] 2.18fF
Xuser_analog_project_wrapper_empty_0 user_analog_project_wrapper_empty_0/gpio_analog[0]
+ user_analog_project_wrapper_empty_0/gpio_analog[10] user_analog_project_wrapper_empty_0/gpio_analog[11]
+ user_analog_project_wrapper_empty_0/gpio_analog[12] user_analog_project_wrapper_empty_0/gpio_analog[13]
+ user_analog_project_wrapper_empty_0/gpio_analog[14] user_analog_project_wrapper_empty_0/gpio_analog[15]
+ user_analog_project_wrapper_empty_0/gpio_analog[16] user_analog_project_wrapper_empty_0/gpio_analog[17]
+ user_analog_project_wrapper_empty_0/gpio_analog[1] user_analog_project_wrapper_empty_0/gpio_analog[2]
+ user_analog_project_wrapper_empty_0/gpio_analog[3] user_analog_project_wrapper_empty_0/gpio_analog[4]
+ user_analog_project_wrapper_empty_0/gpio_analog[5] user_analog_project_wrapper_empty_0/gpio_analog[6]
+ user_analog_project_wrapper_empty_0/gpio_analog[7] user_analog_project_wrapper_empty_0/gpio_analog[8]
+ user_analog_project_wrapper_empty_0/gpio_analog[9] user_analog_project_wrapper_empty_0/gpio_noesd[0]
+ user_analog_project_wrapper_empty_0/gpio_noesd[10] user_analog_project_wrapper_empty_0/gpio_noesd[11]
+ user_analog_project_wrapper_empty_0/gpio_noesd[12] user_analog_project_wrapper_empty_0/gpio_noesd[13]
+ user_analog_project_wrapper_empty_0/gpio_noesd[14] user_analog_project_wrapper_empty_0/gpio_noesd[15]
+ user_analog_project_wrapper_empty_0/gpio_noesd[16] user_analog_project_wrapper_empty_0/gpio_noesd[17]
+ user_analog_project_wrapper_empty_0/gpio_noesd[1] user_analog_project_wrapper_empty_0/gpio_noesd[2]
+ user_analog_project_wrapper_empty_0/gpio_noesd[3] user_analog_project_wrapper_empty_0/gpio_noesd[4]
+ user_analog_project_wrapper_empty_0/gpio_noesd[5] user_analog_project_wrapper_empty_0/gpio_noesd[6]
+ user_analog_project_wrapper_empty_0/gpio_noesd[7] user_analog_project_wrapper_empty_0/gpio_noesd[8]
+ user_analog_project_wrapper_empty_0/gpio_noesd[9] user_analog_project_wrapper_empty_0/io_analog[0]
+ user_analog_project_wrapper_empty_0/io_analog[10] user_analog_project_wrapper_empty_0/io_analog[1]
+ user_analog_project_wrapper_empty_0/io_analog[2] user_analog_project_wrapper_empty_0/io_analog[3]
+ user_analog_project_wrapper_empty_0/io_analog[7] user_analog_project_wrapper_empty_0/io_analog[8]
+ user_analog_project_wrapper_empty_0/io_analog[9] user_analog_project_wrapper_empty_0/io_analog[4]
+ user_analog_project_wrapper_empty_0/io_analog[5] user_analog_project_wrapper_empty_0/io_analog[6]
+ user_analog_project_wrapper_empty_0/io_clamp_high[0] user_analog_project_wrapper_empty_0/io_clamp_high[1]
+ user_analog_project_wrapper_empty_0/io_clamp_high[2] user_analog_project_wrapper_empty_0/io_clamp_low[0]
+ user_analog_project_wrapper_empty_0/io_clamp_low[1] user_analog_project_wrapper_empty_0/io_clamp_low[2]
+ user_analog_project_wrapper_empty_0/io_in[0] user_analog_project_wrapper_empty_0/io_in[10]
+ user_analog_project_wrapper_empty_0/io_in[11] user_analog_project_wrapper_empty_0/io_in[12]
+ user_analog_project_wrapper_empty_0/io_in[13] user_analog_project_wrapper_empty_0/io_in[14]
+ user_analog_project_wrapper_empty_0/io_in[15] user_analog_project_wrapper_empty_0/io_in[16]
+ user_analog_project_wrapper_empty_0/io_in[17] user_analog_project_wrapper_empty_0/io_in[18]
+ user_analog_project_wrapper_empty_0/io_in[19] user_analog_project_wrapper_empty_0/io_in[1]
+ user_analog_project_wrapper_empty_0/io_in[20] user_analog_project_wrapper_empty_0/io_in[21]
+ user_analog_project_wrapper_empty_0/io_in[22] user_analog_project_wrapper_empty_0/io_in[23]
+ user_analog_project_wrapper_empty_0/io_in[24] user_analog_project_wrapper_empty_0/io_in[25]
+ user_analog_project_wrapper_empty_0/io_in[26] user_analog_project_wrapper_empty_0/io_in[2]
+ user_analog_project_wrapper_empty_0/io_in[3] user_analog_project_wrapper_empty_0/io_in[4]
+ user_analog_project_wrapper_empty_0/io_in[5] user_analog_project_wrapper_empty_0/io_in[6]
+ user_analog_project_wrapper_empty_0/io_in[7] user_analog_project_wrapper_empty_0/io_in[8]
+ user_analog_project_wrapper_empty_0/io_in[9] user_analog_project_wrapper_empty_0/io_in_3v3[0]
+ user_analog_project_wrapper_empty_0/io_in_3v3[10] user_analog_project_wrapper_empty_0/io_in_3v3[11]
+ user_analog_project_wrapper_empty_0/io_in_3v3[12] user_analog_project_wrapper_empty_0/io_in_3v3[13]
+ user_analog_project_wrapper_empty_0/io_in_3v3[14] user_analog_project_wrapper_empty_0/io_in_3v3[15]
+ user_analog_project_wrapper_empty_0/io_in_3v3[16] user_analog_project_wrapper_empty_0/io_in_3v3[17]
+ user_analog_project_wrapper_empty_0/io_in_3v3[18] user_analog_project_wrapper_empty_0/io_in_3v3[19]
+ user_analog_project_wrapper_empty_0/io_in_3v3[1] user_analog_project_wrapper_empty_0/io_in_3v3[20]
+ user_analog_project_wrapper_empty_0/io_in_3v3[21] user_analog_project_wrapper_empty_0/io_in_3v3[22]
+ user_analog_project_wrapper_empty_0/io_in_3v3[23] user_analog_project_wrapper_empty_0/io_in_3v3[24]
+ user_analog_project_wrapper_empty_0/io_in_3v3[25] user_analog_project_wrapper_empty_0/io_in_3v3[26]
+ user_analog_project_wrapper_empty_0/io_in_3v3[2] user_analog_project_wrapper_empty_0/io_in_3v3[3]
+ user_analog_project_wrapper_empty_0/io_in_3v3[4] user_analog_project_wrapper_empty_0/io_in_3v3[5]
+ user_analog_project_wrapper_empty_0/io_in_3v3[6] user_analog_project_wrapper_empty_0/io_in_3v3[7]
+ user_analog_project_wrapper_empty_0/io_in_3v3[8] user_analog_project_wrapper_empty_0/io_in_3v3[9]
+ user_analog_project_wrapper_empty_0/io_oeb[0] user_analog_project_wrapper_empty_0/io_oeb[10]
+ user_analog_project_wrapper_empty_0/io_oeb[11] user_analog_project_wrapper_empty_0/io_oeb[12]
+ user_analog_project_wrapper_empty_0/io_oeb[13] user_analog_project_wrapper_empty_0/io_oeb[14]
+ user_analog_project_wrapper_empty_0/io_oeb[15] user_analog_project_wrapper_empty_0/io_oeb[16]
+ user_analog_project_wrapper_empty_0/io_oeb[17] user_analog_project_wrapper_empty_0/io_oeb[18]
+ user_analog_project_wrapper_empty_0/io_oeb[19] user_analog_project_wrapper_empty_0/io_oeb[1]
+ user_analog_project_wrapper_empty_0/io_oeb[20] user_analog_project_wrapper_empty_0/io_oeb[21]
+ user_analog_project_wrapper_empty_0/io_oeb[22] user_analog_project_wrapper_empty_0/io_oeb[23]
+ user_analog_project_wrapper_empty_0/io_oeb[24] user_analog_project_wrapper_empty_0/io_oeb[25]
+ user_analog_project_wrapper_empty_0/io_oeb[26] user_analog_project_wrapper_empty_0/io_oeb[2]
+ user_analog_project_wrapper_empty_0/io_oeb[3] user_analog_project_wrapper_empty_0/io_oeb[4]
+ user_analog_project_wrapper_empty_0/io_oeb[5] user_analog_project_wrapper_empty_0/io_oeb[6]
+ user_analog_project_wrapper_empty_0/io_oeb[7] user_analog_project_wrapper_empty_0/io_oeb[8]
+ user_analog_project_wrapper_empty_0/io_oeb[9] user_analog_project_wrapper_empty_0/io_out[0]
+ user_analog_project_wrapper_empty_0/io_out[10] user_analog_project_wrapper_empty_0/io_out[11]
+ user_analog_project_wrapper_empty_0/io_out[12] user_analog_project_wrapper_empty_0/io_out[13]
+ user_analog_project_wrapper_empty_0/io_out[14] user_analog_project_wrapper_empty_0/io_out[15]
+ user_analog_project_wrapper_empty_0/io_out[16] user_analog_project_wrapper_empty_0/io_out[17]
+ user_analog_project_wrapper_empty_0/io_out[18] user_analog_project_wrapper_empty_0/io_out[19]
+ user_analog_project_wrapper_empty_0/io_out[1] user_analog_project_wrapper_empty_0/io_out[20]
+ user_analog_project_wrapper_empty_0/io_out[21] user_analog_project_wrapper_empty_0/io_out[22]
+ user_analog_project_wrapper_empty_0/io_out[23] user_analog_project_wrapper_empty_0/io_out[24]
+ user_analog_project_wrapper_empty_0/io_out[25] user_analog_project_wrapper_empty_0/io_out[26]
+ user_analog_project_wrapper_empty_0/io_out[2] user_analog_project_wrapper_empty_0/io_out[3]
+ user_analog_project_wrapper_empty_0/io_out[4] user_analog_project_wrapper_empty_0/io_out[5]
+ user_analog_project_wrapper_empty_0/io_out[6] user_analog_project_wrapper_empty_0/io_out[7]
+ user_analog_project_wrapper_empty_0/io_out[8] user_analog_project_wrapper_empty_0/io_out[9]
+ user_analog_project_wrapper_empty_0/la_data_in[0] user_analog_project_wrapper_empty_0/la_data_in[100]
+ user_analog_project_wrapper_empty_0/la_data_in[101] user_analog_project_wrapper_empty_0/la_data_in[102]
+ user_analog_project_wrapper_empty_0/la_data_in[103] user_analog_project_wrapper_empty_0/la_data_in[104]
+ user_analog_project_wrapper_empty_0/la_data_in[105] user_analog_project_wrapper_empty_0/la_data_in[106]
+ user_analog_project_wrapper_empty_0/la_data_in[107] user_analog_project_wrapper_empty_0/la_data_in[108]
+ user_analog_project_wrapper_empty_0/la_data_in[109] user_analog_project_wrapper_empty_0/la_data_in[10]
+ user_analog_project_wrapper_empty_0/la_data_in[110] user_analog_project_wrapper_empty_0/la_data_in[111]
+ user_analog_project_wrapper_empty_0/la_data_in[112] user_analog_project_wrapper_empty_0/la_data_in[113]
+ user_analog_project_wrapper_empty_0/la_data_in[114] user_analog_project_wrapper_empty_0/la_data_in[115]
+ user_analog_project_wrapper_empty_0/la_data_in[116] user_analog_project_wrapper_empty_0/la_data_in[117]
+ user_analog_project_wrapper_empty_0/la_data_in[118] user_analog_project_wrapper_empty_0/la_data_in[119]
+ user_analog_project_wrapper_empty_0/la_data_in[11] user_analog_project_wrapper_empty_0/la_data_in[120]
+ user_analog_project_wrapper_empty_0/la_data_in[121] user_analog_project_wrapper_empty_0/la_data_in[122]
+ user_analog_project_wrapper_empty_0/la_data_in[123] user_analog_project_wrapper_empty_0/la_data_in[124]
+ user_analog_project_wrapper_empty_0/la_data_in[125] user_analog_project_wrapper_empty_0/la_data_in[126]
+ user_analog_project_wrapper_empty_0/la_data_in[127] user_analog_project_wrapper_empty_0/la_data_in[12]
+ user_analog_project_wrapper_empty_0/la_data_in[13] user_analog_project_wrapper_empty_0/la_data_in[14]
+ user_analog_project_wrapper_empty_0/la_data_in[15] user_analog_project_wrapper_empty_0/la_data_in[16]
+ user_analog_project_wrapper_empty_0/la_data_in[17] user_analog_project_wrapper_empty_0/la_data_in[18]
+ user_analog_project_wrapper_empty_0/la_data_in[19] user_analog_project_wrapper_empty_0/la_data_in[1]
+ user_analog_project_wrapper_empty_0/la_data_in[20] user_analog_project_wrapper_empty_0/la_data_in[21]
+ user_analog_project_wrapper_empty_0/la_data_in[22] user_analog_project_wrapper_empty_0/la_data_in[23]
+ user_analog_project_wrapper_empty_0/la_data_in[24] user_analog_project_wrapper_empty_0/la_data_in[25]
+ user_analog_project_wrapper_empty_0/la_data_in[26] user_analog_project_wrapper_empty_0/la_data_in[27]
+ user_analog_project_wrapper_empty_0/la_data_in[28] user_analog_project_wrapper_empty_0/la_data_in[29]
+ user_analog_project_wrapper_empty_0/la_data_in[2] user_analog_project_wrapper_empty_0/la_data_in[30]
+ user_analog_project_wrapper_empty_0/la_data_in[31] user_analog_project_wrapper_empty_0/la_data_in[32]
+ user_analog_project_wrapper_empty_0/la_data_in[33] user_analog_project_wrapper_empty_0/la_data_in[34]
+ user_analog_project_wrapper_empty_0/la_data_in[35] user_analog_project_wrapper_empty_0/la_data_in[36]
+ user_analog_project_wrapper_empty_0/la_data_in[37] user_analog_project_wrapper_empty_0/la_data_in[38]
+ user_analog_project_wrapper_empty_0/la_data_in[39] user_analog_project_wrapper_empty_0/la_data_in[3]
+ user_analog_project_wrapper_empty_0/la_data_in[40] user_analog_project_wrapper_empty_0/la_data_in[41]
+ user_analog_project_wrapper_empty_0/la_data_in[42] user_analog_project_wrapper_empty_0/la_data_in[43]
+ user_analog_project_wrapper_empty_0/la_data_in[44] user_analog_project_wrapper_empty_0/la_data_in[45]
+ user_analog_project_wrapper_empty_0/la_data_in[46] user_analog_project_wrapper_empty_0/la_data_in[47]
+ user_analog_project_wrapper_empty_0/la_data_in[48] user_analog_project_wrapper_empty_0/la_data_in[49]
+ user_analog_project_wrapper_empty_0/la_data_in[4] user_analog_project_wrapper_empty_0/la_data_in[50]
+ user_analog_project_wrapper_empty_0/la_data_in[51] user_analog_project_wrapper_empty_0/la_data_in[52]
+ user_analog_project_wrapper_empty_0/la_data_in[53] user_analog_project_wrapper_empty_0/la_data_in[54]
+ user_analog_project_wrapper_empty_0/la_data_in[55] user_analog_project_wrapper_empty_0/la_data_in[56]
+ user_analog_project_wrapper_empty_0/la_data_in[57] user_analog_project_wrapper_empty_0/la_data_in[58]
+ user_analog_project_wrapper_empty_0/la_data_in[59] user_analog_project_wrapper_empty_0/la_data_in[5]
+ user_analog_project_wrapper_empty_0/la_data_in[60] user_analog_project_wrapper_empty_0/la_data_in[61]
+ user_analog_project_wrapper_empty_0/la_data_in[62] user_analog_project_wrapper_empty_0/la_data_in[63]
+ user_analog_project_wrapper_empty_0/la_data_in[64] user_analog_project_wrapper_empty_0/la_data_in[65]
+ user_analog_project_wrapper_empty_0/la_data_in[66] user_analog_project_wrapper_empty_0/la_data_in[67]
+ user_analog_project_wrapper_empty_0/la_data_in[68] user_analog_project_wrapper_empty_0/la_data_in[69]
+ user_analog_project_wrapper_empty_0/la_data_in[6] user_analog_project_wrapper_empty_0/la_data_in[70]
+ user_analog_project_wrapper_empty_0/la_data_in[71] user_analog_project_wrapper_empty_0/la_data_in[72]
+ user_analog_project_wrapper_empty_0/la_data_in[73] user_analog_project_wrapper_empty_0/la_data_in[74]
+ user_analog_project_wrapper_empty_0/la_data_in[75] user_analog_project_wrapper_empty_0/la_data_in[76]
+ user_analog_project_wrapper_empty_0/la_data_in[77] user_analog_project_wrapper_empty_0/la_data_in[78]
+ user_analog_project_wrapper_empty_0/la_data_in[79] user_analog_project_wrapper_empty_0/la_data_in[7]
+ user_analog_project_wrapper_empty_0/la_data_in[80] user_analog_project_wrapper_empty_0/la_data_in[81]
+ user_analog_project_wrapper_empty_0/la_data_in[82] user_analog_project_wrapper_empty_0/la_data_in[83]
+ user_analog_project_wrapper_empty_0/la_data_in[84] user_analog_project_wrapper_empty_0/la_data_in[85]
+ user_analog_project_wrapper_empty_0/la_data_in[86] user_analog_project_wrapper_empty_0/la_data_in[87]
+ user_analog_project_wrapper_empty_0/la_data_in[88] user_analog_project_wrapper_empty_0/la_data_in[89]
+ user_analog_project_wrapper_empty_0/la_data_in[8] user_analog_project_wrapper_empty_0/la_data_in[90]
+ user_analog_project_wrapper_empty_0/la_data_in[91] user_analog_project_wrapper_empty_0/la_data_in[92]
+ user_analog_project_wrapper_empty_0/la_data_in[93] user_analog_project_wrapper_empty_0/la_data_in[94]
+ user_analog_project_wrapper_empty_0/la_data_in[95] user_analog_project_wrapper_empty_0/la_data_in[96]
+ user_analog_project_wrapper_empty_0/la_data_in[97] user_analog_project_wrapper_empty_0/la_data_in[98]
+ user_analog_project_wrapper_empty_0/la_data_in[99] user_analog_project_wrapper_empty_0/la_data_in[9]
+ user_analog_project_wrapper_empty_0/la_data_out[0] user_analog_project_wrapper_empty_0/la_data_out[100]
+ user_analog_project_wrapper_empty_0/la_data_out[101] user_analog_project_wrapper_empty_0/la_data_out[102]
+ user_analog_project_wrapper_empty_0/la_data_out[103] user_analog_project_wrapper_empty_0/la_data_out[104]
+ user_analog_project_wrapper_empty_0/la_data_out[105] user_analog_project_wrapper_empty_0/la_data_out[106]
+ user_analog_project_wrapper_empty_0/la_data_out[107] user_analog_project_wrapper_empty_0/la_data_out[108]
+ user_analog_project_wrapper_empty_0/la_data_out[109] user_analog_project_wrapper_empty_0/la_data_out[10]
+ user_analog_project_wrapper_empty_0/la_data_out[110] user_analog_project_wrapper_empty_0/la_data_out[111]
+ user_analog_project_wrapper_empty_0/la_data_out[112] user_analog_project_wrapper_empty_0/la_data_out[113]
+ user_analog_project_wrapper_empty_0/la_data_out[114] user_analog_project_wrapper_empty_0/la_data_out[115]
+ user_analog_project_wrapper_empty_0/la_data_out[116] user_analog_project_wrapper_empty_0/la_data_out[117]
+ user_analog_project_wrapper_empty_0/la_data_out[118] user_analog_project_wrapper_empty_0/la_data_out[119]
+ user_analog_project_wrapper_empty_0/la_data_out[11] user_analog_project_wrapper_empty_0/la_data_out[120]
+ user_analog_project_wrapper_empty_0/la_data_out[121] user_analog_project_wrapper_empty_0/la_data_out[122]
+ user_analog_project_wrapper_empty_0/la_data_out[123] user_analog_project_wrapper_empty_0/la_data_out[124]
+ user_analog_project_wrapper_empty_0/la_data_out[125] user_analog_project_wrapper_empty_0/la_data_out[126]
+ user_analog_project_wrapper_empty_0/la_data_out[127] user_analog_project_wrapper_empty_0/la_data_out[12]
+ user_analog_project_wrapper_empty_0/la_data_out[13] user_analog_project_wrapper_empty_0/la_data_out[14]
+ user_analog_project_wrapper_empty_0/la_data_out[15] user_analog_project_wrapper_empty_0/la_data_out[16]
+ user_analog_project_wrapper_empty_0/la_data_out[17] user_analog_project_wrapper_empty_0/la_data_out[18]
+ user_analog_project_wrapper_empty_0/la_data_out[19] user_analog_project_wrapper_empty_0/la_data_out[1]
+ user_analog_project_wrapper_empty_0/la_data_out[20] user_analog_project_wrapper_empty_0/la_data_out[21]
+ user_analog_project_wrapper_empty_0/la_data_out[22] user_analog_project_wrapper_empty_0/la_data_out[23]
+ user_analog_project_wrapper_empty_0/la_data_out[24] user_analog_project_wrapper_empty_0/la_data_out[25]
+ user_analog_project_wrapper_empty_0/la_data_out[26] user_analog_project_wrapper_empty_0/la_data_out[27]
+ user_analog_project_wrapper_empty_0/la_data_out[28] user_analog_project_wrapper_empty_0/la_data_out[29]
+ user_analog_project_wrapper_empty_0/la_data_out[2] user_analog_project_wrapper_empty_0/la_data_out[30]
+ user_analog_project_wrapper_empty_0/la_data_out[31] user_analog_project_wrapper_empty_0/la_data_out[32]
+ user_analog_project_wrapper_empty_0/la_data_out[33] user_analog_project_wrapper_empty_0/la_data_out[34]
+ user_analog_project_wrapper_empty_0/la_data_out[35] user_analog_project_wrapper_empty_0/la_data_out[36]
+ user_analog_project_wrapper_empty_0/la_data_out[37] user_analog_project_wrapper_empty_0/la_data_out[38]
+ user_analog_project_wrapper_empty_0/la_data_out[39] user_analog_project_wrapper_empty_0/la_data_out[3]
+ user_analog_project_wrapper_empty_0/la_data_out[40] user_analog_project_wrapper_empty_0/la_data_out[41]
+ user_analog_project_wrapper_empty_0/la_data_out[42] user_analog_project_wrapper_empty_0/la_data_out[43]
+ user_analog_project_wrapper_empty_0/la_data_out[44] user_analog_project_wrapper_empty_0/la_data_out[45]
+ user_analog_project_wrapper_empty_0/la_data_out[46] user_analog_project_wrapper_empty_0/la_data_out[47]
+ user_analog_project_wrapper_empty_0/la_data_out[48] user_analog_project_wrapper_empty_0/la_data_out[49]
+ user_analog_project_wrapper_empty_0/la_data_out[4] user_analog_project_wrapper_empty_0/la_data_out[50]
+ user_analog_project_wrapper_empty_0/la_data_out[51] user_analog_project_wrapper_empty_0/la_data_out[52]
+ user_analog_project_wrapper_empty_0/la_data_out[53] user_analog_project_wrapper_empty_0/la_data_out[54]
+ user_analog_project_wrapper_empty_0/la_data_out[55] user_analog_project_wrapper_empty_0/la_data_out[56]
+ user_analog_project_wrapper_empty_0/la_data_out[57] user_analog_project_wrapper_empty_0/la_data_out[58]
+ user_analog_project_wrapper_empty_0/la_data_out[59] user_analog_project_wrapper_empty_0/la_data_out[5]
+ user_analog_project_wrapper_empty_0/la_data_out[60] user_analog_project_wrapper_empty_0/la_data_out[61]
+ user_analog_project_wrapper_empty_0/la_data_out[62] user_analog_project_wrapper_empty_0/la_data_out[63]
+ user_analog_project_wrapper_empty_0/la_data_out[64] user_analog_project_wrapper_empty_0/la_data_out[65]
+ user_analog_project_wrapper_empty_0/la_data_out[66] user_analog_project_wrapper_empty_0/la_data_out[67]
+ user_analog_project_wrapper_empty_0/la_data_out[68] user_analog_project_wrapper_empty_0/la_data_out[69]
+ user_analog_project_wrapper_empty_0/la_data_out[6] user_analog_project_wrapper_empty_0/la_data_out[70]
+ user_analog_project_wrapper_empty_0/la_data_out[71] user_analog_project_wrapper_empty_0/la_data_out[72]
+ user_analog_project_wrapper_empty_0/la_data_out[73] user_analog_project_wrapper_empty_0/la_data_out[74]
+ user_analog_project_wrapper_empty_0/la_data_out[75] user_analog_project_wrapper_empty_0/la_data_out[76]
+ user_analog_project_wrapper_empty_0/la_data_out[77] user_analog_project_wrapper_empty_0/la_data_out[78]
+ user_analog_project_wrapper_empty_0/la_data_out[79] user_analog_project_wrapper_empty_0/la_data_out[7]
+ user_analog_project_wrapper_empty_0/la_data_out[80] user_analog_project_wrapper_empty_0/la_data_out[81]
+ user_analog_project_wrapper_empty_0/la_data_out[82] user_analog_project_wrapper_empty_0/la_data_out[83]
+ user_analog_project_wrapper_empty_0/la_data_out[84] user_analog_project_wrapper_empty_0/la_data_out[85]
+ user_analog_project_wrapper_empty_0/la_data_out[86] user_analog_project_wrapper_empty_0/la_data_out[87]
+ user_analog_project_wrapper_empty_0/la_data_out[88] user_analog_project_wrapper_empty_0/la_data_out[89]
+ user_analog_project_wrapper_empty_0/la_data_out[8] user_analog_project_wrapper_empty_0/la_data_out[90]
+ user_analog_project_wrapper_empty_0/la_data_out[91] user_analog_project_wrapper_empty_0/la_data_out[92]
+ user_analog_project_wrapper_empty_0/la_data_out[93] user_analog_project_wrapper_empty_0/la_data_out[94]
+ user_analog_project_wrapper_empty_0/la_data_out[95] user_analog_project_wrapper_empty_0/la_data_out[96]
+ user_analog_project_wrapper_empty_0/la_data_out[97] user_analog_project_wrapper_empty_0/la_data_out[98]
+ user_analog_project_wrapper_empty_0/la_data_out[99] user_analog_project_wrapper_empty_0/la_data_out[9]
+ user_analog_project_wrapper_empty_0/la_oenb[0] user_analog_project_wrapper_empty_0/la_oenb[100]
+ user_analog_project_wrapper_empty_0/la_oenb[101] user_analog_project_wrapper_empty_0/la_oenb[102]
+ user_analog_project_wrapper_empty_0/la_oenb[103] user_analog_project_wrapper_empty_0/la_oenb[104]
+ user_analog_project_wrapper_empty_0/la_oenb[105] user_analog_project_wrapper_empty_0/la_oenb[106]
+ user_analog_project_wrapper_empty_0/la_oenb[107] user_analog_project_wrapper_empty_0/la_oenb[108]
+ user_analog_project_wrapper_empty_0/la_oenb[109] user_analog_project_wrapper_empty_0/la_oenb[10]
+ user_analog_project_wrapper_empty_0/la_oenb[110] user_analog_project_wrapper_empty_0/la_oenb[111]
+ user_analog_project_wrapper_empty_0/la_oenb[112] user_analog_project_wrapper_empty_0/la_oenb[113]
+ user_analog_project_wrapper_empty_0/la_oenb[114] user_analog_project_wrapper_empty_0/la_oenb[115]
+ user_analog_project_wrapper_empty_0/la_oenb[116] user_analog_project_wrapper_empty_0/la_oenb[117]
+ user_analog_project_wrapper_empty_0/la_oenb[118] user_analog_project_wrapper_empty_0/la_oenb[119]
+ user_analog_project_wrapper_empty_0/la_oenb[11] user_analog_project_wrapper_empty_0/la_oenb[120]
+ user_analog_project_wrapper_empty_0/la_oenb[121] user_analog_project_wrapper_empty_0/la_oenb[122]
+ user_analog_project_wrapper_empty_0/la_oenb[123] user_analog_project_wrapper_empty_0/la_oenb[124]
+ user_analog_project_wrapper_empty_0/la_oenb[125] user_analog_project_wrapper_empty_0/la_oenb[126]
+ user_analog_project_wrapper_empty_0/la_oenb[127] user_analog_project_wrapper_empty_0/la_oenb[12]
+ user_analog_project_wrapper_empty_0/la_oenb[13] user_analog_project_wrapper_empty_0/la_oenb[14]
+ user_analog_project_wrapper_empty_0/la_oenb[15] user_analog_project_wrapper_empty_0/la_oenb[16]
+ user_analog_project_wrapper_empty_0/la_oenb[17] user_analog_project_wrapper_empty_0/la_oenb[18]
+ user_analog_project_wrapper_empty_0/la_oenb[19] user_analog_project_wrapper_empty_0/la_oenb[1]
+ user_analog_project_wrapper_empty_0/la_oenb[20] user_analog_project_wrapper_empty_0/la_oenb[21]
+ user_analog_project_wrapper_empty_0/la_oenb[22] user_analog_project_wrapper_empty_0/la_oenb[23]
+ user_analog_project_wrapper_empty_0/la_oenb[24] user_analog_project_wrapper_empty_0/la_oenb[25]
+ user_analog_project_wrapper_empty_0/la_oenb[26] user_analog_project_wrapper_empty_0/la_oenb[27]
+ user_analog_project_wrapper_empty_0/la_oenb[28] user_analog_project_wrapper_empty_0/la_oenb[29]
+ user_analog_project_wrapper_empty_0/la_oenb[2] user_analog_project_wrapper_empty_0/la_oenb[30]
+ user_analog_project_wrapper_empty_0/la_oenb[31] user_analog_project_wrapper_empty_0/la_oenb[32]
+ user_analog_project_wrapper_empty_0/la_oenb[33] user_analog_project_wrapper_empty_0/la_oenb[34]
+ user_analog_project_wrapper_empty_0/la_oenb[35] user_analog_project_wrapper_empty_0/la_oenb[36]
+ user_analog_project_wrapper_empty_0/la_oenb[37] user_analog_project_wrapper_empty_0/la_oenb[38]
+ user_analog_project_wrapper_empty_0/la_oenb[39] user_analog_project_wrapper_empty_0/la_oenb[3]
+ user_analog_project_wrapper_empty_0/la_oenb[40] user_analog_project_wrapper_empty_0/la_oenb[41]
+ user_analog_project_wrapper_empty_0/la_oenb[42] user_analog_project_wrapper_empty_0/la_oenb[43]
+ user_analog_project_wrapper_empty_0/la_oenb[44] user_analog_project_wrapper_empty_0/la_oenb[45]
+ user_analog_project_wrapper_empty_0/la_oenb[46] user_analog_project_wrapper_empty_0/la_oenb[47]
+ user_analog_project_wrapper_empty_0/la_oenb[48] user_analog_project_wrapper_empty_0/la_oenb[49]
+ user_analog_project_wrapper_empty_0/la_oenb[4] user_analog_project_wrapper_empty_0/la_oenb[50]
+ user_analog_project_wrapper_empty_0/la_oenb[51] user_analog_project_wrapper_empty_0/la_oenb[52]
+ user_analog_project_wrapper_empty_0/la_oenb[53] user_analog_project_wrapper_empty_0/la_oenb[54]
+ user_analog_project_wrapper_empty_0/la_oenb[55] user_analog_project_wrapper_empty_0/la_oenb[56]
+ user_analog_project_wrapper_empty_0/la_oenb[57] user_analog_project_wrapper_empty_0/la_oenb[58]
+ user_analog_project_wrapper_empty_0/la_oenb[59] user_analog_project_wrapper_empty_0/la_oenb[5]
+ user_analog_project_wrapper_empty_0/la_oenb[60] user_analog_project_wrapper_empty_0/la_oenb[61]
+ user_analog_project_wrapper_empty_0/la_oenb[62] user_analog_project_wrapper_empty_0/la_oenb[63]
+ user_analog_project_wrapper_empty_0/la_oenb[64] user_analog_project_wrapper_empty_0/la_oenb[65]
+ user_analog_project_wrapper_empty_0/la_oenb[66] user_analog_project_wrapper_empty_0/la_oenb[67]
+ user_analog_project_wrapper_empty_0/la_oenb[68] user_analog_project_wrapper_empty_0/la_oenb[69]
+ user_analog_project_wrapper_empty_0/la_oenb[6] user_analog_project_wrapper_empty_0/la_oenb[70]
+ user_analog_project_wrapper_empty_0/la_oenb[71] user_analog_project_wrapper_empty_0/la_oenb[72]
+ user_analog_project_wrapper_empty_0/la_oenb[73] user_analog_project_wrapper_empty_0/la_oenb[74]
+ user_analog_project_wrapper_empty_0/la_oenb[75] user_analog_project_wrapper_empty_0/la_oenb[76]
+ user_analog_project_wrapper_empty_0/la_oenb[77] user_analog_project_wrapper_empty_0/la_oenb[78]
+ user_analog_project_wrapper_empty_0/la_oenb[79] user_analog_project_wrapper_empty_0/la_oenb[7]
+ user_analog_project_wrapper_empty_0/la_oenb[80] user_analog_project_wrapper_empty_0/la_oenb[81]
+ user_analog_project_wrapper_empty_0/la_oenb[82] user_analog_project_wrapper_empty_0/la_oenb[83]
+ user_analog_project_wrapper_empty_0/la_oenb[84] user_analog_project_wrapper_empty_0/la_oenb[85]
+ user_analog_project_wrapper_empty_0/la_oenb[86] user_analog_project_wrapper_empty_0/la_oenb[87]
+ user_analog_project_wrapper_empty_0/la_oenb[88] user_analog_project_wrapper_empty_0/la_oenb[89]
+ user_analog_project_wrapper_empty_0/la_oenb[8] user_analog_project_wrapper_empty_0/la_oenb[90]
+ user_analog_project_wrapper_empty_0/la_oenb[91] user_analog_project_wrapper_empty_0/la_oenb[92]
+ user_analog_project_wrapper_empty_0/la_oenb[93] user_analog_project_wrapper_empty_0/la_oenb[94]
+ user_analog_project_wrapper_empty_0/la_oenb[95] user_analog_project_wrapper_empty_0/la_oenb[96]
+ user_analog_project_wrapper_empty_0/la_oenb[97] user_analog_project_wrapper_empty_0/la_oenb[98]
+ user_analog_project_wrapper_empty_0/la_oenb[99] user_analog_project_wrapper_empty_0/la_oenb[9]
+ user_analog_project_wrapper_empty_0/user_clock2 user_analog_project_wrapper_empty_0/user_irq[0]
+ user_analog_project_wrapper_empty_0/user_irq[1] user_analog_project_wrapper_empty_0/user_irq[2]
+ user_analog_project_wrapper_empty_0/vccd1 user_analog_project_wrapper_empty_0/vccd2
+ user_analog_project_wrapper_empty_0/vdda1 user_analog_project_wrapper_empty_0/vdda2
+ VSUBS user_analog_project_wrapper_empty_0/vssa2 user_analog_project_wrapper_empty_0/vssd1
+ user_analog_project_wrapper_empty_0/vssd2 user_analog_project_wrapper_empty_0/wb_clk_i
+ user_analog_project_wrapper_empty_0/wb_rst_i user_analog_project_wrapper_empty_0/wbs_ack_o
+ user_analog_project_wrapper_empty_0/wbs_adr_i[0] user_analog_project_wrapper_empty_0/wbs_adr_i[10]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[11] user_analog_project_wrapper_empty_0/wbs_adr_i[12]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[13] user_analog_project_wrapper_empty_0/wbs_adr_i[14]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[15] user_analog_project_wrapper_empty_0/wbs_adr_i[16]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[17] user_analog_project_wrapper_empty_0/wbs_adr_i[18]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[19] user_analog_project_wrapper_empty_0/wbs_adr_i[1]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[20] user_analog_project_wrapper_empty_0/wbs_adr_i[21]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[22] user_analog_project_wrapper_empty_0/wbs_adr_i[23]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[24] user_analog_project_wrapper_empty_0/wbs_adr_i[25]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[26] user_analog_project_wrapper_empty_0/wbs_adr_i[27]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[28] user_analog_project_wrapper_empty_0/wbs_adr_i[29]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[2] user_analog_project_wrapper_empty_0/wbs_adr_i[30]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[31] user_analog_project_wrapper_empty_0/wbs_adr_i[3]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[4] user_analog_project_wrapper_empty_0/wbs_adr_i[5]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[6] user_analog_project_wrapper_empty_0/wbs_adr_i[7]
+ user_analog_project_wrapper_empty_0/wbs_adr_i[8] user_analog_project_wrapper_empty_0/wbs_adr_i[9]
+ user_analog_project_wrapper_empty_0/wbs_cyc_i user_analog_project_wrapper_empty_0/wbs_dat_i[0]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[10] user_analog_project_wrapper_empty_0/wbs_dat_i[11]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[12] user_analog_project_wrapper_empty_0/wbs_dat_i[13]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[14] user_analog_project_wrapper_empty_0/wbs_dat_i[15]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[16] user_analog_project_wrapper_empty_0/wbs_dat_i[17]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[18] user_analog_project_wrapper_empty_0/wbs_dat_i[19]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[1] user_analog_project_wrapper_empty_0/wbs_dat_i[20]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[21] user_analog_project_wrapper_empty_0/wbs_dat_i[22]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[23] user_analog_project_wrapper_empty_0/wbs_dat_i[24]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[25] user_analog_project_wrapper_empty_0/wbs_dat_i[26]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[27] user_analog_project_wrapper_empty_0/wbs_dat_i[28]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[29] user_analog_project_wrapper_empty_0/wbs_dat_i[2]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[30] user_analog_project_wrapper_empty_0/wbs_dat_i[31]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[3] user_analog_project_wrapper_empty_0/wbs_dat_i[4]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[5] user_analog_project_wrapper_empty_0/wbs_dat_i[6]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[7] user_analog_project_wrapper_empty_0/wbs_dat_i[8]
+ user_analog_project_wrapper_empty_0/wbs_dat_i[9] user_analog_project_wrapper_empty_0/wbs_dat_o[0]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[10] user_analog_project_wrapper_empty_0/wbs_dat_o[11]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[12] user_analog_project_wrapper_empty_0/wbs_dat_o[13]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[14] user_analog_project_wrapper_empty_0/wbs_dat_o[15]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[16] user_analog_project_wrapper_empty_0/wbs_dat_o[17]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[18] user_analog_project_wrapper_empty_0/wbs_dat_o[19]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[1] user_analog_project_wrapper_empty_0/wbs_dat_o[20]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[21] user_analog_project_wrapper_empty_0/wbs_dat_o[22]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[23] user_analog_project_wrapper_empty_0/wbs_dat_o[24]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[25] user_analog_project_wrapper_empty_0/wbs_dat_o[26]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[27] user_analog_project_wrapper_empty_0/wbs_dat_o[28]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[29] user_analog_project_wrapper_empty_0/wbs_dat_o[2]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[30] user_analog_project_wrapper_empty_0/wbs_dat_o[31]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[3] user_analog_project_wrapper_empty_0/wbs_dat_o[4]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[5] user_analog_project_wrapper_empty_0/wbs_dat_o[6]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[7] user_analog_project_wrapper_empty_0/wbs_dat_o[8]
+ user_analog_project_wrapper_empty_0/wbs_dat_o[9] user_analog_project_wrapper_empty_0/wbs_sel_i[0]
+ user_analog_project_wrapper_empty_0/wbs_sel_i[1] user_analog_project_wrapper_empty_0/wbs_sel_i[2]
+ user_analog_project_wrapper_empty_0/wbs_sel_i[3] user_analog_project_wrapper_empty_0/wbs_stb_i
+ user_analog_project_wrapper_empty_0/wbs_we_i user_analog_project_wrapper_empty
Xuser_analog_proj_example_0/ulqc_ldo_0 user_analog_project_wrapper_empty_0/io_analog[0]
+ user_analog_project_wrapper_empty_0/io_analog[4] user_analog_project_wrapper_empty_0/io_analog[5]
+ user_analog_project_wrapper_empty_0/io_analog[6] VSUBS user_analog_project_wrapper_empty_0/io_analog[7]
+ user_analog_project_wrapper_empty_0/vssa2 user_analog_project_wrapper_empty_0/vssd1
+ user_analog_project_wrapper_empty_0/io_analog[8] user_analog_project_wrapper_empty_0/io_analog[1]
+ user_analog_project_wrapper_empty_0/io_analog[9] user_analog_proj_example_0/ulqc_ldo_0/VIN2
+ user_analog_project_wrapper_empty_0/io_analog[10] user_analog_project_wrapper_empty_0/vdda2
+ ulqc_ldo
Xulqc_ldo_0 ulqc_ldo_0/ADJ ulqc_ldo_0/BGRT1 ulqc_ldo_0/BGRT2 ulqc_ldo_0/BGR_OUT VSUBS
+ ulqc_ldo_0/EA_OUT ulqc_ldo_0/VSS2 ulqc_ldo_0/VSS3 ulqc_ldo_0/VOUT1 ulqc_ldo_0/VIN1
+ ulqc_ldo_0/VOUT2 ulqc_ldo_0/VIN2 ulqc_ldo_0/VOUT3 ulqc_ldo_0/VIN3 ulqc_ldo
C16 user_analog_project_wrapper_empty_0/io_analog[7] VSUBS 244.90fF
C17 user_analog_project_wrapper_empty_0/vdda2 VSUBS 641.68fF
C18 user_analog_project_wrapper_empty_0/vssd1 VSUBS 502.55fF
C19 user_analog_project_wrapper_empty_0/io_analog[10] VSUBS 564.58fF
C20 user_analog_proj_example_0/ulqc_ldo_0/VIN2 VSUBS 24.86fF
C21 user_analog_project_wrapper_empty_0/io_analog[9] VSUBS 258.86fF
C22 user_analog_project_wrapper_empty_0/vssa2 VSUBS 346.26fF
C23 user_analog_project_wrapper_empty_0/io_analog[0] VSUBS 328.95fF
C24 user_analog_project_wrapper_empty_0/io_analog[4] VSUBS 226.56fF
C25 user_analog_project_wrapper_empty_0/io_analog[1] VSUBS 143.65fF
C26 user_analog_project_wrapper_empty_0/io_analog[8] VSUBS 420.23fF
C27 user_analog_project_wrapper_empty_0/io_analog[5] VSUBS 158.86fF
C28 user_analog_project_wrapper_empty_0/io_analog[6] VSUBS 326.18fF
C29 user_analog_project_wrapper_empty_0/vssd2 VSUBS 13.26fF
C30 user_analog_project_wrapper_empty_0/vdda1 VSUBS 26.51fF
C31 user_analog_project_wrapper_empty_0/vccd1 VSUBS 13.26fF
C32 user_analog_project_wrapper_empty_0/vccd2 VSUBS 13.26fF
C33 user_analog_project_wrapper_empty_0/io_analog[2] VSUBS 6.94fF
C34 user_analog_project_wrapper_empty_0/io_analog[3] VSUBS 6.94fF
C35 user_analog_project_wrapper_empty_0/io_clamp_high[0] VSUBS 2.83fF
C36 user_analog_project_wrapper_empty_0/io_clamp_low[0] VSUBS 2.83fF
C37 user_analog_project_wrapper_empty_0/io_clamp_high[1] VSUBS 2.83fF
C38 user_analog_project_wrapper_empty_0/io_clamp_low[1] VSUBS 2.83fF
C39 user_analog_project_wrapper_empty_0/io_clamp_high[2] VSUBS 2.83fF
C40 user_analog_project_wrapper_empty_0/io_clamp_low[2] VSUBS 2.83fF
