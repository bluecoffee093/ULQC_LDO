magic
tech sky130A
magscale 1 2
timestamp 1698059623
<< error_p >>
rect -796 581 -738 587
rect -678 581 -620 587
rect -560 581 -502 587
rect -442 581 -384 587
rect -324 581 -266 587
rect -206 581 -148 587
rect -88 581 -30 587
rect 30 581 88 587
rect 148 581 206 587
rect 266 581 324 587
rect 384 581 442 587
rect 502 581 560 587
rect 620 581 678 587
rect 738 581 796 587
rect -796 547 -784 581
rect -678 547 -666 581
rect -560 547 -548 581
rect -442 547 -430 581
rect -324 547 -312 581
rect -206 547 -194 581
rect -88 547 -76 581
rect 30 547 42 581
rect 148 547 160 581
rect 266 547 278 581
rect 384 547 396 581
rect 502 547 514 581
rect 620 547 632 581
rect 738 547 750 581
rect -796 541 -738 547
rect -678 541 -620 547
rect -560 541 -502 547
rect -442 541 -384 547
rect -324 541 -266 547
rect -206 541 -148 547
rect -88 541 -30 547
rect 30 541 88 547
rect 148 541 206 547
rect 266 541 324 547
rect 384 541 442 547
rect 502 541 560 547
rect 620 541 678 547
rect 738 541 796 547
rect -796 -547 -738 -541
rect -678 -547 -620 -541
rect -560 -547 -502 -541
rect -442 -547 -384 -541
rect -324 -547 -266 -541
rect -206 -547 -148 -541
rect -88 -547 -30 -541
rect 30 -547 88 -541
rect 148 -547 206 -541
rect 266 -547 324 -541
rect 384 -547 442 -541
rect 502 -547 560 -541
rect 620 -547 678 -541
rect 738 -547 796 -541
rect -796 -581 -784 -547
rect -678 -581 -666 -547
rect -560 -581 -548 -547
rect -442 -581 -430 -547
rect -324 -581 -312 -547
rect -206 -581 -194 -547
rect -88 -581 -76 -547
rect 30 -581 42 -547
rect 148 -581 160 -547
rect 266 -581 278 -547
rect 384 -581 396 -547
rect 502 -581 514 -547
rect 620 -581 632 -547
rect 738 -581 750 -547
rect -796 -587 -738 -581
rect -678 -587 -620 -581
rect -560 -587 -502 -581
rect -442 -587 -384 -581
rect -324 -587 -266 -581
rect -206 -587 -148 -581
rect -88 -587 -30 -581
rect 30 -587 88 -581
rect 148 -587 206 -581
rect 266 -587 324 -581
rect 384 -587 442 -581
rect 502 -587 560 -581
rect 620 -587 678 -581
rect 738 -587 796 -581
<< nwell >>
rect -993 -719 993 719
<< pmos >>
rect -797 -500 -737 500
rect -679 -500 -619 500
rect -561 -500 -501 500
rect -443 -500 -383 500
rect -325 -500 -265 500
rect -207 -500 -147 500
rect -89 -500 -29 500
rect 29 -500 89 500
rect 147 -500 207 500
rect 265 -500 325 500
rect 383 -500 443 500
rect 501 -500 561 500
rect 619 -500 679 500
rect 737 -500 797 500
<< pdiff >>
rect -855 488 -797 500
rect -855 -488 -843 488
rect -809 -488 -797 488
rect -855 -500 -797 -488
rect -737 488 -679 500
rect -737 -488 -725 488
rect -691 -488 -679 488
rect -737 -500 -679 -488
rect -619 488 -561 500
rect -619 -488 -607 488
rect -573 -488 -561 488
rect -619 -500 -561 -488
rect -501 488 -443 500
rect -501 -488 -489 488
rect -455 -488 -443 488
rect -501 -500 -443 -488
rect -383 488 -325 500
rect -383 -488 -371 488
rect -337 -488 -325 488
rect -383 -500 -325 -488
rect -265 488 -207 500
rect -265 -488 -253 488
rect -219 -488 -207 488
rect -265 -500 -207 -488
rect -147 488 -89 500
rect -147 -488 -135 488
rect -101 -488 -89 488
rect -147 -500 -89 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 89 488 147 500
rect 89 -488 101 488
rect 135 -488 147 488
rect 89 -500 147 -488
rect 207 488 265 500
rect 207 -488 219 488
rect 253 -488 265 488
rect 207 -500 265 -488
rect 325 488 383 500
rect 325 -488 337 488
rect 371 -488 383 488
rect 325 -500 383 -488
rect 443 488 501 500
rect 443 -488 455 488
rect 489 -488 501 488
rect 443 -500 501 -488
rect 561 488 619 500
rect 561 -488 573 488
rect 607 -488 619 488
rect 561 -500 619 -488
rect 679 488 737 500
rect 679 -488 691 488
rect 725 -488 737 488
rect 679 -500 737 -488
rect 797 488 855 500
rect 797 -488 809 488
rect 843 -488 855 488
rect 797 -500 855 -488
<< pdiffc >>
rect -843 -488 -809 488
rect -725 -488 -691 488
rect -607 -488 -573 488
rect -489 -488 -455 488
rect -371 -488 -337 488
rect -253 -488 -219 488
rect -135 -488 -101 488
rect -17 -488 17 488
rect 101 -488 135 488
rect 219 -488 253 488
rect 337 -488 371 488
rect 455 -488 489 488
rect 573 -488 607 488
rect 691 -488 725 488
rect 809 -488 843 488
<< nsubdiff >>
rect -957 649 -861 683
rect 861 649 957 683
rect -957 587 -923 649
rect 923 587 957 649
rect -957 -649 -923 -587
rect 923 -649 957 -587
rect -957 -683 -861 -649
rect 861 -683 957 -649
<< nsubdiffcont >>
rect -861 649 861 683
rect -957 -587 -923 587
rect 923 -587 957 587
rect -861 -683 861 -649
<< poly >>
rect -800 581 -734 597
rect -800 547 -784 581
rect -750 547 -734 581
rect -800 531 -734 547
rect -682 581 -616 597
rect -682 547 -666 581
rect -632 547 -616 581
rect -682 531 -616 547
rect -564 581 -498 597
rect -564 547 -548 581
rect -514 547 -498 581
rect -564 531 -498 547
rect -446 581 -380 597
rect -446 547 -430 581
rect -396 547 -380 581
rect -446 531 -380 547
rect -328 581 -262 597
rect -328 547 -312 581
rect -278 547 -262 581
rect -328 531 -262 547
rect -210 581 -144 597
rect -210 547 -194 581
rect -160 547 -144 581
rect -210 531 -144 547
rect -92 581 -26 597
rect -92 547 -76 581
rect -42 547 -26 581
rect -92 531 -26 547
rect 26 581 92 597
rect 26 547 42 581
rect 76 547 92 581
rect 26 531 92 547
rect 144 581 210 597
rect 144 547 160 581
rect 194 547 210 581
rect 144 531 210 547
rect 262 581 328 597
rect 262 547 278 581
rect 312 547 328 581
rect 262 531 328 547
rect 380 581 446 597
rect 380 547 396 581
rect 430 547 446 581
rect 380 531 446 547
rect 498 581 564 597
rect 498 547 514 581
rect 548 547 564 581
rect 498 531 564 547
rect 616 581 682 597
rect 616 547 632 581
rect 666 547 682 581
rect 616 531 682 547
rect 734 581 800 597
rect 734 547 750 581
rect 784 547 800 581
rect 734 531 800 547
rect -797 500 -737 531
rect -679 500 -619 531
rect -561 500 -501 531
rect -443 500 -383 531
rect -325 500 -265 531
rect -207 500 -147 531
rect -89 500 -29 531
rect 29 500 89 531
rect 147 500 207 531
rect 265 500 325 531
rect 383 500 443 531
rect 501 500 561 531
rect 619 500 679 531
rect 737 500 797 531
rect -797 -531 -737 -500
rect -679 -531 -619 -500
rect -561 -531 -501 -500
rect -443 -531 -383 -500
rect -325 -531 -265 -500
rect -207 -531 -147 -500
rect -89 -531 -29 -500
rect 29 -531 89 -500
rect 147 -531 207 -500
rect 265 -531 325 -500
rect 383 -531 443 -500
rect 501 -531 561 -500
rect 619 -531 679 -500
rect 737 -531 797 -500
rect -800 -547 -734 -531
rect -800 -581 -784 -547
rect -750 -581 -734 -547
rect -800 -597 -734 -581
rect -682 -547 -616 -531
rect -682 -581 -666 -547
rect -632 -581 -616 -547
rect -682 -597 -616 -581
rect -564 -547 -498 -531
rect -564 -581 -548 -547
rect -514 -581 -498 -547
rect -564 -597 -498 -581
rect -446 -547 -380 -531
rect -446 -581 -430 -547
rect -396 -581 -380 -547
rect -446 -597 -380 -581
rect -328 -547 -262 -531
rect -328 -581 -312 -547
rect -278 -581 -262 -547
rect -328 -597 -262 -581
rect -210 -547 -144 -531
rect -210 -581 -194 -547
rect -160 -581 -144 -547
rect -210 -597 -144 -581
rect -92 -547 -26 -531
rect -92 -581 -76 -547
rect -42 -581 -26 -547
rect -92 -597 -26 -581
rect 26 -547 92 -531
rect 26 -581 42 -547
rect 76 -581 92 -547
rect 26 -597 92 -581
rect 144 -547 210 -531
rect 144 -581 160 -547
rect 194 -581 210 -547
rect 144 -597 210 -581
rect 262 -547 328 -531
rect 262 -581 278 -547
rect 312 -581 328 -547
rect 262 -597 328 -581
rect 380 -547 446 -531
rect 380 -581 396 -547
rect 430 -581 446 -547
rect 380 -597 446 -581
rect 498 -547 564 -531
rect 498 -581 514 -547
rect 548 -581 564 -547
rect 498 -597 564 -581
rect 616 -547 682 -531
rect 616 -581 632 -547
rect 666 -581 682 -547
rect 616 -597 682 -581
rect 734 -547 800 -531
rect 734 -581 750 -547
rect 784 -581 800 -547
rect 734 -597 800 -581
<< polycont >>
rect -784 547 -750 581
rect -666 547 -632 581
rect -548 547 -514 581
rect -430 547 -396 581
rect -312 547 -278 581
rect -194 547 -160 581
rect -76 547 -42 581
rect 42 547 76 581
rect 160 547 194 581
rect 278 547 312 581
rect 396 547 430 581
rect 514 547 548 581
rect 632 547 666 581
rect 750 547 784 581
rect -784 -581 -750 -547
rect -666 -581 -632 -547
rect -548 -581 -514 -547
rect -430 -581 -396 -547
rect -312 -581 -278 -547
rect -194 -581 -160 -547
rect -76 -581 -42 -547
rect 42 -581 76 -547
rect 160 -581 194 -547
rect 278 -581 312 -547
rect 396 -581 430 -547
rect 514 -581 548 -547
rect 632 -581 666 -547
rect 750 -581 784 -547
<< locali >>
rect -957 649 -861 683
rect 861 649 957 683
rect -957 587 -923 649
rect 923 587 957 649
rect -800 547 -784 581
rect -750 547 -734 581
rect -682 547 -666 581
rect -632 547 -616 581
rect -564 547 -548 581
rect -514 547 -498 581
rect -446 547 -430 581
rect -396 547 -380 581
rect -328 547 -312 581
rect -278 547 -262 581
rect -210 547 -194 581
rect -160 547 -144 581
rect -92 547 -76 581
rect -42 547 -26 581
rect 26 547 42 581
rect 76 547 92 581
rect 144 547 160 581
rect 194 547 210 581
rect 262 547 278 581
rect 312 547 328 581
rect 380 547 396 581
rect 430 547 446 581
rect 498 547 514 581
rect 548 547 564 581
rect 616 547 632 581
rect 666 547 682 581
rect 734 547 750 581
rect 784 547 800 581
rect -843 488 -809 504
rect -843 -504 -809 -488
rect -725 488 -691 504
rect -725 -504 -691 -488
rect -607 488 -573 504
rect -607 -504 -573 -488
rect -489 488 -455 504
rect -489 -504 -455 -488
rect -371 488 -337 504
rect -371 -504 -337 -488
rect -253 488 -219 504
rect -253 -504 -219 -488
rect -135 488 -101 504
rect -135 -504 -101 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 101 488 135 504
rect 101 -504 135 -488
rect 219 488 253 504
rect 219 -504 253 -488
rect 337 488 371 504
rect 337 -504 371 -488
rect 455 488 489 504
rect 455 -504 489 -488
rect 573 488 607 504
rect 573 -504 607 -488
rect 691 488 725 504
rect 691 -504 725 -488
rect 809 488 843 504
rect 809 -504 843 -488
rect -800 -581 -784 -547
rect -750 -581 -734 -547
rect -682 -581 -666 -547
rect -632 -581 -616 -547
rect -564 -581 -548 -547
rect -514 -581 -498 -547
rect -446 -581 -430 -547
rect -396 -581 -380 -547
rect -328 -581 -312 -547
rect -278 -581 -262 -547
rect -210 -581 -194 -547
rect -160 -581 -144 -547
rect -92 -581 -76 -547
rect -42 -581 -26 -547
rect 26 -581 42 -547
rect 76 -581 92 -547
rect 144 -581 160 -547
rect 194 -581 210 -547
rect 262 -581 278 -547
rect 312 -581 328 -547
rect 380 -581 396 -547
rect 430 -581 446 -547
rect 498 -581 514 -547
rect 548 -581 564 -547
rect 616 -581 632 -547
rect 666 -581 682 -547
rect 734 -581 750 -547
rect 784 -581 800 -547
rect -957 -649 -923 -587
rect 923 -649 957 -587
rect -957 -683 -861 -649
rect 861 -683 957 -649
<< viali >>
rect -784 547 -750 581
rect -666 547 -632 581
rect -548 547 -514 581
rect -430 547 -396 581
rect -312 547 -278 581
rect -194 547 -160 581
rect -76 547 -42 581
rect 42 547 76 581
rect 160 547 194 581
rect 278 547 312 581
rect 396 547 430 581
rect 514 547 548 581
rect 632 547 666 581
rect 750 547 784 581
rect -843 -488 -809 488
rect -725 -488 -691 488
rect -607 -488 -573 488
rect -489 -488 -455 488
rect -371 -488 -337 488
rect -253 -488 -219 488
rect -135 -488 -101 488
rect -17 -488 17 488
rect 101 -488 135 488
rect 219 -488 253 488
rect 337 -488 371 488
rect 455 -488 489 488
rect 573 -488 607 488
rect 691 -488 725 488
rect 809 -488 843 488
rect -784 -581 -750 -547
rect -666 -581 -632 -547
rect -548 -581 -514 -547
rect -430 -581 -396 -547
rect -312 -581 -278 -547
rect -194 -581 -160 -547
rect -76 -581 -42 -547
rect 42 -581 76 -547
rect 160 -581 194 -547
rect 278 -581 312 -547
rect 396 -581 430 -547
rect 514 -581 548 -547
rect 632 -581 666 -547
rect 750 -581 784 -547
<< metal1 >>
rect -796 581 -738 587
rect -796 547 -784 581
rect -750 547 -738 581
rect -796 541 -738 547
rect -678 581 -620 587
rect -678 547 -666 581
rect -632 547 -620 581
rect -678 541 -620 547
rect -560 581 -502 587
rect -560 547 -548 581
rect -514 547 -502 581
rect -560 541 -502 547
rect -442 581 -384 587
rect -442 547 -430 581
rect -396 547 -384 581
rect -442 541 -384 547
rect -324 581 -266 587
rect -324 547 -312 581
rect -278 547 -266 581
rect -324 541 -266 547
rect -206 581 -148 587
rect -206 547 -194 581
rect -160 547 -148 581
rect -206 541 -148 547
rect -88 581 -30 587
rect -88 547 -76 581
rect -42 547 -30 581
rect -88 541 -30 547
rect 30 581 88 587
rect 30 547 42 581
rect 76 547 88 581
rect 30 541 88 547
rect 148 581 206 587
rect 148 547 160 581
rect 194 547 206 581
rect 148 541 206 547
rect 266 581 324 587
rect 266 547 278 581
rect 312 547 324 581
rect 266 541 324 547
rect 384 581 442 587
rect 384 547 396 581
rect 430 547 442 581
rect 384 541 442 547
rect 502 581 560 587
rect 502 547 514 581
rect 548 547 560 581
rect 502 541 560 547
rect 620 581 678 587
rect 620 547 632 581
rect 666 547 678 581
rect 620 541 678 547
rect 738 581 796 587
rect 738 547 750 581
rect 784 547 796 581
rect 738 541 796 547
rect -849 488 -803 500
rect -849 -488 -843 488
rect -809 -488 -803 488
rect -849 -500 -803 -488
rect -731 488 -685 500
rect -731 -488 -725 488
rect -691 -488 -685 488
rect -731 -500 -685 -488
rect -613 488 -567 500
rect -613 -488 -607 488
rect -573 -488 -567 488
rect -613 -500 -567 -488
rect -495 488 -449 500
rect -495 -488 -489 488
rect -455 -488 -449 488
rect -495 -500 -449 -488
rect -377 488 -331 500
rect -377 -488 -371 488
rect -337 -488 -331 488
rect -377 -500 -331 -488
rect -259 488 -213 500
rect -259 -488 -253 488
rect -219 -488 -213 488
rect -259 -500 -213 -488
rect -141 488 -95 500
rect -141 -488 -135 488
rect -101 -488 -95 488
rect -141 -500 -95 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 95 488 141 500
rect 95 -488 101 488
rect 135 -488 141 488
rect 95 -500 141 -488
rect 213 488 259 500
rect 213 -488 219 488
rect 253 -488 259 488
rect 213 -500 259 -488
rect 331 488 377 500
rect 331 -488 337 488
rect 371 -488 377 488
rect 331 -500 377 -488
rect 449 488 495 500
rect 449 -488 455 488
rect 489 -488 495 488
rect 449 -500 495 -488
rect 567 488 613 500
rect 567 -488 573 488
rect 607 -488 613 488
rect 567 -500 613 -488
rect 685 488 731 500
rect 685 -488 691 488
rect 725 -488 731 488
rect 685 -500 731 -488
rect 803 488 849 500
rect 803 -488 809 488
rect 843 -488 849 488
rect 803 -500 849 -488
rect -796 -547 -738 -541
rect -796 -581 -784 -547
rect -750 -581 -738 -547
rect -796 -587 -738 -581
rect -678 -547 -620 -541
rect -678 -581 -666 -547
rect -632 -581 -620 -547
rect -678 -587 -620 -581
rect -560 -547 -502 -541
rect -560 -581 -548 -547
rect -514 -581 -502 -547
rect -560 -587 -502 -581
rect -442 -547 -384 -541
rect -442 -581 -430 -547
rect -396 -581 -384 -547
rect -442 -587 -384 -581
rect -324 -547 -266 -541
rect -324 -581 -312 -547
rect -278 -581 -266 -547
rect -324 -587 -266 -581
rect -206 -547 -148 -541
rect -206 -581 -194 -547
rect -160 -581 -148 -547
rect -206 -587 -148 -581
rect -88 -547 -30 -541
rect -88 -581 -76 -547
rect -42 -581 -30 -547
rect -88 -587 -30 -581
rect 30 -547 88 -541
rect 30 -581 42 -547
rect 76 -581 88 -547
rect 30 -587 88 -581
rect 148 -547 206 -541
rect 148 -581 160 -547
rect 194 -581 206 -547
rect 148 -587 206 -581
rect 266 -547 324 -541
rect 266 -581 278 -547
rect 312 -581 324 -547
rect 266 -587 324 -581
rect 384 -547 442 -541
rect 384 -581 396 -547
rect 430 -581 442 -547
rect 384 -587 442 -581
rect 502 -547 560 -541
rect 502 -581 514 -547
rect 548 -581 560 -547
rect 502 -587 560 -581
rect 620 -547 678 -541
rect 620 -581 632 -547
rect 666 -581 678 -547
rect 620 -587 678 -581
rect 738 -547 796 -541
rect 738 -581 750 -547
rect 784 -581 796 -547
rect 738 -587 796 -581
<< properties >>
string FIXED_BBOX -940 -666 940 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 0.3 m 1 nf 14 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
