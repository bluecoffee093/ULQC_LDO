magic
tech sky130A
magscale 1 2
timestamp 1695677300
<< metal1 >>
rect 249328 588174 249586 593942
rect 249328 587972 250806 588174
rect 247854 587464 250470 587664
rect 250948 587466 251148 592642
rect 251292 587940 251532 592000
rect 252198 587900 252438 591960
rect 250594 587096 250604 587296
rect 250804 587096 250814 587296
rect 251266 587096 251276 587296
rect 251476 587096 251486 587296
rect 251846 587086 251856 587286
rect 252056 587086 252066 587286
rect 252462 587084 252472 587284
rect 252672 587084 252682 587284
rect 252910 587092 253892 587290
rect 248284 586712 250438 586912
rect 248530 586276 250684 586476
rect 250958 585256 251176 586904
rect 253028 586276 255986 586490
<< via1 >>
rect 250604 587096 250804 587296
rect 251276 587096 251476 587296
rect 251856 587086 252056 587286
rect 252472 587084 252672 587284
<< metal2 >>
rect 250604 587296 250804 587306
rect 246604 587096 250604 587296
rect 250604 587086 250804 587096
rect 251276 587296 251476 587306
rect 251276 585488 251476 587096
rect 251856 587286 252056 587296
rect 251856 585362 252056 587086
rect 252472 587284 252672 587294
rect 252472 585100 252672 587084
use user_analog_proj_example  user_analog_proj_example_0
timestamp 1695673762
transform 1 0 245230 0 1 578608
box 5008 7668 7940 9565
use user_analog_project_wrapper_empty  user_analog_project_wrapper_empty_0
timestamp 1632839657
transform 1 0 0 0 1 0
box -800 -800 584800 704800
<< end >>
