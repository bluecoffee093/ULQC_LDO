magic
tech sky130A
magscale 1 2
timestamp 1696967143
<< checkpaint >>
rect -1366 99791 3546 99844
rect -1366 99685 5885 99791
rect -1366 -766 10563 99685
rect 973 -819 10563 -766
rect 3312 -872 10563 -819
rect 5651 -925 10563 -872
use sky130_fd_pr__pfet_01v8_lvt_B5ZT88  XM1
timestamp 0
transform 1 0 1090 0 1 49539
box -1196 -49045 1196 49045
use sky130_fd_pr__pfet_01v8_lvt_B5ZT88  XM2
timestamp 0
transform 1 0 3429 0 1 49486
box -1196 -49045 1196 49045
use sky130_fd_pr__nfet_01v8_2DGCRD  XM3
timestamp 0
transform 1 0 5768 0 1 49361
box -1196 -48973 1196 48973
use sky130_fd_pr__nfet_01v8_2DGCRD  XM4
timestamp 0
transform 1 0 1143 0 1 49520
box -1196 -48973 1196 48973
use sky130_fd_pr__pfet_01v8_lvt_B5ZT88  XM5
timestamp 0
transform 1 0 8107 0 1 49380
box -1196 -49045 1196 49045
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1675710598
transform 1 0 2339 0 1 547
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ2
array 0 0 796 0 7 796
timestamp 1675710598
transform 1 0 -53 0 1 547
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ3
timestamp 1675710598
transform 1 0 3135 0 1 547
box 0 0 796 796
<< end >>
