* NGSPICE file created from power_transistor.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_KPD88M w_n785_n300# a_15_n200# a_n561_n200# a_n177_n200#
+ a_111_n200# a_n129_n297# a_n513_n297# a_n609_231# a_n273_n200# a_63_n297# a_n749_n200#
+ a_687_n200# a_n321_n297# a_159_231# a_639_n297# a_n81_n200# a_399_n200# a_351_231#
+ a_495_n200# a_n33_231# a_447_n297# a_n225_231# a_591_n200# a_n657_n200# a_207_n200#
+ a_543_231# a_n369_n200# a_303_n200# a_n705_n297# a_255_n297# a_n417_231# a_n465_n200#
X0 a_n657_n200# a_n705_n297# a_n749_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X1 a_n273_n200# a_n321_n297# a_n369_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_303_n200# a_255_n297# a_207_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_591_n200# a_543_231# a_495_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_n177_n200# a_n225_231# a_n273_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X5 a_207_n200# a_159_231# a_111_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_495_n200# a_447_n297# a_399_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_n561_n200# a_n609_231# a_n657_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X8 a_111_n200# a_63_n297# a_15_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X9 a_399_n200# a_351_231# a_303_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 a_n465_n200# a_n513_n297# a_n561_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X11 a_687_n200# a_639_n297# a_591_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X12 a_n81_n200# a_n129_n297# a_n177_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X13 a_15_n200# a_n33_231# a_n81_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 a_n369_n200# a_n417_231# a_n465_n200# w_n785_n300# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt power_transistor VDD EA_OUT OUT BIAS_CURR
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|0] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|1] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|2] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|3] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|4] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|5] VDD BIAS_CURR BIAS_CURR BIAS_CURR VDD EA_OUT
+ EA_OUT EA_OUT VDD EA_OUT BIAS_CURR VDD EA_OUT EA_OUT EA_OUT VDD BIAS_CURR EA_OUT
+ VDD EA_OUT EA_OUT EA_OUT BIAS_CURR VDD BIAS_CURR EA_OUT BIAS_CURR VDD EA_OUT EA_OUT
+ EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|5] VDD BIAS_CURR BIAS_CURR BIAS_CURR VDD EA_OUT
+ EA_OUT EA_OUT VDD EA_OUT BIAS_CURR VDD EA_OUT EA_OUT EA_OUT VDD BIAS_CURR EA_OUT
+ VDD EA_OUT EA_OUT EA_OUT BIAS_CURR VDD BIAS_CURR EA_OUT BIAS_CURR VDD EA_OUT EA_OUT
+ EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|5] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|6] VDD BIAS_CURR BIAS_CURR BIAS_CURR VDD EA_OUT
+ EA_OUT EA_OUT VDD EA_OUT BIAS_CURR VDD EA_OUT EA_OUT EA_OUT VDD BIAS_CURR EA_OUT
+ VDD EA_OUT EA_OUT EA_OUT BIAS_CURR VDD BIAS_CURR EA_OUT BIAS_CURR VDD EA_OUT EA_OUT
+ EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|6] VDD BIAS_CURR BIAS_CURR BIAS_CURR VDD EA_OUT
+ EA_OUT EA_OUT VDD EA_OUT BIAS_CURR VDD EA_OUT EA_OUT EA_OUT VDD BIAS_CURR EA_OUT
+ VDD EA_OUT EA_OUT EA_OUT BIAS_CURR VDD BIAS_CURR EA_OUT BIAS_CURR VDD EA_OUT EA_OUT
+ EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|6] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|7] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|8] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|9] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|10] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[0|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[1|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[2|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[3|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[4|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[5|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[6|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[7|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[8|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[9|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD
+ EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT OUT
+ VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[10|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[11|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[12|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[13|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[14|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[15|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[16|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[17|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[18|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[19|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[20|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[21|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[22|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[23|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[24|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[25|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[26|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[27|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[28|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
Xsky130_fd_pr__pfet_01v8_KPD88M_0[29|11] VDD OUT OUT OUT VDD EA_OUT EA_OUT EA_OUT
+ VDD EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD OUT EA_OUT VDD EA_OUT EA_OUT EA_OUT
+ OUT VDD OUT EA_OUT OUT VDD EA_OUT EA_OUT EA_OUT VDD sky130_fd_pr__pfet_01v8_KPD88M
*R0 OUT m3_9940_11524# sky130_fd_pr__res_generic_m3 w=3.55e+06u l=50000u
*R1 VDD m3_10968_9535# sky130_fd_pr__res_generic_m3 w=3.55e+06u l=50000u
*R2 OUT m3_11768_11524# sky130_fd_pr__res_generic_m3 w=3.55e+06u l=50000u
*R3 VDD m3_9140_9535# sky130_fd_pr__res_generic_m3 w=3.55e+06u l=50000u
.ends

