magic
tech sky130A
magscale 1 2
timestamp 1697794495
<< error_p >>
rect -88 545 -30 551
rect 30 545 88 551
rect -88 511 -76 545
rect 30 511 42 545
rect -88 505 -30 511
rect 30 505 88 511
<< nwell >>
rect -183 -598 183 564
<< pmos >>
rect -89 -536 -29 464
rect 29 -536 89 464
<< pdiff >>
rect -147 452 -89 464
rect -147 -524 -135 452
rect -101 -524 -89 452
rect -147 -536 -89 -524
rect -29 452 29 464
rect -29 -524 -17 452
rect 17 -524 29 452
rect -29 -536 29 -524
rect 89 452 147 464
rect 89 -524 101 452
rect 135 -524 147 452
rect 89 -536 147 -524
<< pdiffc >>
rect -135 -524 -101 452
rect -17 -524 17 452
rect 101 -524 135 452
<< poly >>
rect -92 545 -26 561
rect -92 511 -76 545
rect -42 511 -26 545
rect -92 495 -26 511
rect 26 545 92 561
rect 26 511 42 545
rect 76 511 92 545
rect 26 495 92 511
rect -89 464 -29 495
rect 29 464 89 495
rect -89 -562 -29 -536
rect 29 -562 89 -536
<< polycont >>
rect -76 511 -42 545
rect 42 511 76 545
<< locali >>
rect -92 511 -76 545
rect -42 511 -26 545
rect 26 511 42 545
rect 76 511 92 545
rect -135 452 -101 468
rect -135 -540 -101 -524
rect -17 452 17 468
rect -17 -540 17 -524
rect 101 452 135 468
rect 101 -540 135 -524
<< viali >>
rect -76 511 -42 545
rect 42 511 76 545
rect -135 -524 -101 452
rect -17 -524 17 452
rect 101 -524 135 452
<< metal1 >>
rect -88 545 -30 551
rect -88 511 -76 545
rect -42 511 -30 545
rect -88 505 -30 511
rect 30 545 88 551
rect 30 511 42 545
rect 76 511 88 545
rect 30 505 88 511
rect -141 452 -95 464
rect -141 -524 -135 452
rect -101 -524 -95 452
rect -141 -536 -95 -524
rect -23 452 23 464
rect -23 -524 -17 452
rect 17 -524 23 452
rect -23 -536 23 -524
rect 95 452 141 464
rect 95 -524 101 452
rect 135 -524 141 452
rect 95 -536 141 -524
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 0.3 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
