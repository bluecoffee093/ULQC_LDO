magic
tech sky130A
magscale 1 2
timestamp 1697796765
<< nwell >>
rect -183 -562 183 562
<< pmos >>
rect -89 -500 -29 500
rect 29 -500 89 500
<< pdiff >>
rect -147 488 -89 500
rect -147 -488 -135 488
rect -101 -488 -89 488
rect -147 -500 -89 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 89 488 147 500
rect 89 -488 101 488
rect 135 -488 147 488
rect 89 -500 147 -488
<< pdiffc >>
rect -135 -488 -101 488
rect -17 -488 17 488
rect 101 -488 135 488
<< poly >>
rect -89 500 -29 526
rect 29 500 89 526
rect -89 -526 -29 -500
rect 29 -526 89 -500
<< locali >>
rect -135 488 -101 504
rect -135 -504 -101 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 101 488 135 504
rect 101 -504 135 -488
<< viali >>
rect -135 -488 -101 488
rect -17 -488 17 488
rect 101 -488 135 488
<< metal1 >>
rect -141 488 -95 500
rect -141 -488 -135 488
rect -101 -488 -95 488
rect -141 -500 -95 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 95 488 141 500
rect 95 -488 101 488
rect 135 -488 141 488
rect 95 -500 141 -488
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 0.3 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
