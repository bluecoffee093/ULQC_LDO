magic
tech sky130A
magscale 1 2
timestamp 1697811681
<< nmos >>
rect -1261 -1000 -1061 1000
rect -1003 -1000 -803 1000
rect -745 -1000 -545 1000
rect -487 -1000 -287 1000
rect -229 -1000 -29 1000
rect 29 -1000 229 1000
rect 287 -1000 487 1000
rect 545 -1000 745 1000
rect 803 -1000 1003 1000
rect 1061 -1000 1261 1000
<< ndiff >>
rect -1319 988 -1261 1000
rect -1319 -988 -1307 988
rect -1273 -988 -1261 988
rect -1319 -1000 -1261 -988
rect -1061 988 -1003 1000
rect -1061 -988 -1049 988
rect -1015 -988 -1003 988
rect -1061 -1000 -1003 -988
rect -803 988 -745 1000
rect -803 -988 -791 988
rect -757 -988 -745 988
rect -803 -1000 -745 -988
rect -545 988 -487 1000
rect -545 -988 -533 988
rect -499 -988 -487 988
rect -545 -1000 -487 -988
rect -287 988 -229 1000
rect -287 -988 -275 988
rect -241 -988 -229 988
rect -287 -1000 -229 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 229 988 287 1000
rect 229 -988 241 988
rect 275 -988 287 988
rect 229 -1000 287 -988
rect 487 988 545 1000
rect 487 -988 499 988
rect 533 -988 545 988
rect 487 -1000 545 -988
rect 745 988 803 1000
rect 745 -988 757 988
rect 791 -988 803 988
rect 745 -1000 803 -988
rect 1003 988 1061 1000
rect 1003 -988 1015 988
rect 1049 -988 1061 988
rect 1003 -1000 1061 -988
rect 1261 988 1319 1000
rect 1261 -988 1273 988
rect 1307 -988 1319 988
rect 1261 -1000 1319 -988
<< ndiffc >>
rect -1307 -988 -1273 988
rect -1049 -988 -1015 988
rect -791 -988 -757 988
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
rect 757 -988 791 988
rect 1015 -988 1049 988
rect 1273 -988 1307 988
<< poly >>
rect -1261 1000 -1061 1026
rect -1003 1000 -803 1026
rect -745 1000 -545 1026
rect -487 1000 -287 1026
rect -229 1000 -29 1026
rect 29 1000 229 1026
rect 287 1000 487 1026
rect 545 1000 745 1026
rect 803 1000 1003 1026
rect 1061 1000 1261 1026
rect -1261 -1026 -1061 -1000
rect -1003 -1026 -803 -1000
rect -745 -1026 -545 -1000
rect -487 -1026 -287 -1000
rect -229 -1026 -29 -1000
rect 29 -1026 229 -1000
rect 287 -1026 487 -1000
rect 545 -1026 745 -1000
rect 803 -1026 1003 -1000
rect 1061 -1026 1261 -1000
<< locali >>
rect -1307 988 -1273 1004
rect -1307 -1004 -1273 -988
rect -1049 988 -1015 1004
rect -1049 -1004 -1015 -988
rect -791 988 -757 1004
rect -791 -1004 -757 -988
rect -533 988 -499 1004
rect -533 -1004 -499 -988
rect -275 988 -241 1004
rect -275 -1004 -241 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 241 988 275 1004
rect 241 -1004 275 -988
rect 499 988 533 1004
rect 499 -1004 533 -988
rect 757 988 791 1004
rect 757 -1004 791 -988
rect 1015 988 1049 1004
rect 1015 -1004 1049 -988
rect 1273 988 1307 1004
rect 1273 -1004 1307 -988
<< viali >>
rect -1307 -988 -1273 988
rect -1049 -988 -1015 988
rect -791 -988 -757 988
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
rect 757 -988 791 988
rect 1015 -988 1049 988
rect 1273 -988 1307 988
<< metal1 >>
rect -1313 988 -1267 1000
rect -1313 -988 -1307 988
rect -1273 -988 -1267 988
rect -1313 -1000 -1267 -988
rect -1055 988 -1009 1000
rect -1055 -988 -1049 988
rect -1015 -988 -1009 988
rect -1055 -1000 -1009 -988
rect -797 988 -751 1000
rect -797 -988 -791 988
rect -757 -988 -751 988
rect -797 -1000 -751 -988
rect -539 988 -493 1000
rect -539 -988 -533 988
rect -499 -988 -493 988
rect -539 -1000 -493 -988
rect -281 988 -235 1000
rect -281 -988 -275 988
rect -241 -988 -235 988
rect -281 -1000 -235 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 235 988 281 1000
rect 235 -988 241 988
rect 275 -988 281 988
rect 235 -1000 281 -988
rect 493 988 539 1000
rect 493 -988 499 988
rect 533 -988 539 988
rect 493 -1000 539 -988
rect 751 988 797 1000
rect 751 -988 757 988
rect 791 -988 797 988
rect 751 -1000 797 -988
rect 1009 988 1055 1000
rect 1009 -988 1015 988
rect 1049 -988 1055 988
rect 1009 -1000 1055 -988
rect 1267 988 1313 1000
rect 1267 -988 1273 988
rect 1307 -988 1313 988
rect 1267 -1000 1313 -988
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 1 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
