magic
tech sky130A
magscale 1 2
timestamp 1698945223
<< metal2 >>
rect 465400 699400 470400 699410
rect 453100 696600 465400 699400
rect 453100 696590 470400 696600
rect 453100 634300 467300 696590
rect 443200 632800 447600 632810
rect 447600 631600 453600 632800
rect 443200 631590 447600 631600
rect 439400 628700 453800 630900
rect 439400 628600 444600 628700
rect 439400 624590 444600 624600
<< via2 >>
rect 465400 696600 470400 699400
rect 443200 631600 447600 632800
rect 439400 624600 444600 628600
<< metal3 >>
rect 120200 628600 125200 704800
rect 413400 698700 418400 704800
rect 465400 699405 470400 704800
rect 465390 699400 470410 699405
rect 413400 695300 447600 698700
rect 465390 696600 465400 699400
rect 470400 696600 470410 699400
rect 465390 696595 470410 696600
rect 443200 632805 447600 695300
rect 510600 694100 525400 704800
rect 510590 686100 510600 694100
rect 525400 686100 525410 694100
rect 572690 666700 572700 683000
rect 580700 678000 584000 683000
rect 580700 666700 580710 678000
rect 443190 632800 447610 632805
rect 443190 631600 443200 632800
rect 447600 631600 447610 632800
rect 443190 631595 447610 631600
rect 439390 628600 444610 628605
rect 120200 624600 439400 628600
rect 444600 624600 444610 628600
rect 439390 624595 444610 624600
<< via3 >>
rect 510600 686100 525400 694100
rect 572700 666700 580700 683000
<< metal4 >>
rect 510599 694100 525401 694101
rect 510599 686100 510600 694100
rect 525400 686100 525401 694100
rect 510599 686099 525401 686100
rect 572699 683000 580701 683001
rect 318450 681598 497270 681600
rect 318450 669082 318996 681598
rect 334292 681594 497270 681598
rect 334292 669082 489270 681594
rect 318450 669078 489270 669082
rect 572699 666700 572700 683000
rect 580700 666700 580701 683000
rect 572699 666699 580701 666700
<< via4 >>
rect 510600 686100 525400 694100
rect 318996 669082 334292 681598
rect 489270 669078 497284 681594
rect 572700 666700 580700 683000
rect 452201 616122 460201 624122
<< metal5 >>
rect 318994 701916 323994 702300
rect 329294 701916 334294 702300
rect 318994 681622 334294 701916
rect 510576 694100 525424 694124
rect 452200 686100 510600 694100
rect 525400 686100 525700 694100
rect 318972 681598 334316 681622
rect 318972 669082 318996 681598
rect 334292 669082 334316 681598
rect 318972 669058 334316 669082
rect 452201 624146 460201 686100
rect 510576 686076 525424 686100
rect 572676 683000 580724 683024
rect 489246 681594 497308 681618
rect 489246 669078 489270 681594
rect 497284 669078 497308 681594
rect 489246 669054 497308 669078
rect 489270 651482 497270 669054
rect 572676 666700 572700 683000
rect 580700 666700 580724 683000
rect 572676 666676 580724 666700
rect 572700 651200 580700 666676
rect 497800 643200 580700 651200
rect 452177 624122 460225 624146
rect 452177 616122 452201 624122
rect 460201 616122 460225 624122
rect 452177 616098 460225 616122
use ulqc_ldo  ulqc_ldo_0
timestamp 1698945223
transform 1 0 455019 0 1 620414
box -2065 -11200 50651 31068
use user_analog_project_wrapper_empty  user_analog_project_wrapper_empty_0
timestamp 1632839657
transform 1 0 0 0 1 0
box -800 -800 584800 704800
<< end >>
