magic
tech sky130A
magscale 1 2
timestamp 1695692044
<< metal1 >>
rect 229234 699750 230288 699890
rect 229234 699376 229326 699750
rect 230220 699376 230288 699750
rect 70042 696412 71614 696752
rect 70042 694638 70200 696412
rect 71346 694638 71614 696412
rect 70042 588912 71614 694638
rect 70014 587298 227256 588912
rect 229234 588054 230288 699376
rect 318996 697144 323898 697254
rect 318996 696784 319098 697144
rect 323672 696784 323898 697144
rect 249330 671696 249588 671700
rect 318996 671696 323898 696784
rect 560904 682638 579550 682990
rect 560904 678578 577306 682638
rect 578930 678578 579550 682638
rect 560904 677982 579550 678578
rect 249330 671354 323898 671696
rect 249330 593942 249588 671354
rect 318996 669538 323898 671354
rect 560946 646680 561550 677982
rect 251288 646316 561550 646680
rect 251288 646312 561548 646316
rect 249328 593844 249588 593942
rect 249328 588174 249586 593844
rect 250940 592422 250950 592644
rect 251150 592422 251160 592644
rect 70014 587150 224660 587298
rect 224650 587146 224660 587150
rect 227262 587146 227272 587298
rect 229238 586488 230284 588054
rect 249328 587972 250806 588174
rect 247854 587662 250470 587664
rect 247848 587460 247858 587662
rect 248062 587464 250470 587662
rect 250948 587466 251148 592422
rect 251290 592000 251530 646312
rect 253596 613054 253606 616202
rect 253900 613054 253910 616202
rect 253604 612158 253906 613054
rect 251290 591866 251532 592000
rect 251292 587940 251532 591866
rect 252188 590848 252198 591564
rect 252436 590848 252446 591564
rect 252198 587900 252438 590848
rect 248062 587460 248072 587464
rect 250594 587096 250604 587296
rect 250804 587096 250814 587296
rect 251266 587096 251276 587296
rect 251476 587096 251486 587296
rect 253618 587290 253898 612158
rect 570052 593918 570062 594480
rect 570460 593918 570470 594480
rect 258596 593592 259018 593620
rect 258586 593088 258596 593592
rect 259020 593088 259030 593592
rect 251846 587086 251856 587286
rect 252056 587086 252066 587286
rect 252462 587084 252472 587284
rect 252672 587084 252682 587284
rect 252910 587092 253898 587290
rect 253618 587086 253898 587092
rect 248284 586910 250438 586912
rect 248282 586712 250438 586910
rect 229230 586474 247574 586488
rect 229230 586274 247246 586474
rect 247576 586274 247586 586474
rect 229230 586256 247574 586274
rect 79356 585498 79366 585500
rect 51584 585254 79366 585498
rect 79672 585254 79682 585500
rect 51584 564244 57966 585254
rect 17818 563802 57978 564244
rect 17818 559876 18390 563802
rect 24696 559876 57978 563802
rect 17818 559410 57978 559876
rect 51584 559372 57966 559410
rect 61492 536482 61502 536716
rect 61792 536712 61802 536716
rect 61792 536694 72312 536712
rect 61792 536484 71970 536694
rect 72312 536484 72322 536694
rect 61792 536482 61802 536484
rect 10326 499348 10336 500976
rect 12198 500952 12208 500976
rect 75784 500952 75794 500954
rect 12198 499350 75794 500952
rect 78128 499350 78138 500954
rect 12198 499348 12208 499350
rect 248282 474848 248542 586712
rect 249000 586472 250684 586476
rect 248994 586274 249004 586472
rect 249250 586276 250684 586472
rect 249250 586274 249260 586276
rect 250958 585502 251176 586904
rect 253744 586490 253986 586492
rect 253028 586276 255986 586490
rect 250948 585256 250958 585502
rect 251176 585256 251186 585502
rect 248278 311944 248544 474848
rect 248272 311796 248544 311944
rect 248272 168786 248538 311796
rect 253744 197748 253986 586276
rect 258596 585284 259018 593088
rect 570062 590196 570462 593918
rect 570058 589920 570068 590196
rect 570462 589920 570472 590196
rect 570062 589918 570462 589920
rect 258588 585090 258598 585284
rect 259018 585090 259028 585284
rect 258596 585088 259018 585090
rect 253744 197546 567938 197748
rect 253744 197538 253986 197546
rect 565856 195368 567938 197546
rect 565856 182656 566304 195368
rect 567232 182656 567938 195368
rect 565856 181418 567938 182656
rect 572374 168800 574026 168816
rect 572072 168798 574026 168800
rect 519508 168786 574026 168798
rect 248268 168380 574026 168786
rect 519508 168374 574026 168380
rect 572374 151048 574026 168374
rect 572374 137846 572678 151048
rect 573596 137846 574026 151048
rect 572374 136838 574026 137846
<< via1 >>
rect 229326 699376 230220 699750
rect 70200 694638 71346 696412
rect 319098 696784 323672 697144
rect 577306 678578 578930 682638
rect 250950 592422 251150 592644
rect 224660 587146 227262 587298
rect 247858 587460 248062 587662
rect 253606 613054 253900 616202
rect 252198 590848 252436 591564
rect 250604 587096 250804 587296
rect 251276 587096 251476 587296
rect 570062 593918 570460 594480
rect 258596 593088 259020 593592
rect 251856 587086 252056 587286
rect 252472 587084 252672 587284
rect 247246 586274 247576 586474
rect 79366 585254 79672 585500
rect 18390 559876 24696 563802
rect 61502 536482 61792 536716
rect 71970 536484 72312 536694
rect 10336 499348 12198 500976
rect 75794 499350 78128 500954
rect 249004 586274 249250 586472
rect 250958 585256 251176 585502
rect 570068 589920 570462 590196
rect 258598 585090 259018 585284
rect 566304 182656 567232 195368
rect 572678 137846 573596 151048
<< metal2 >>
rect 229326 699750 230220 699760
rect 229326 699366 230220 699376
rect 32758 699214 33394 699280
rect 16202 698414 33394 699214
rect 16202 696930 16760 698414
rect 19950 696930 33394 698414
rect 570062 698478 570456 698566
rect 16202 696096 33394 696930
rect 177234 697256 180314 697868
rect 10390 685002 12190 685176
rect 10390 680624 10510 685002
rect 11920 680624 12190 685002
rect 10390 500986 12190 680624
rect 18390 563802 24696 563812
rect 18390 559866 24696 559876
rect 32758 536716 33394 696096
rect 70200 696412 71346 696422
rect 70200 694628 71346 694638
rect 177234 695890 177698 697256
rect 179686 695890 180314 697256
rect 570062 697722 570110 698478
rect 570364 697722 570456 698478
rect 319098 697144 323672 697154
rect 319098 696774 323672 696784
rect 121900 694248 123554 694480
rect 121900 692996 122082 694248
rect 123324 692996 123554 694248
rect 121900 594118 123554 692996
rect 177234 616562 180314 695890
rect 570062 657162 570456 697722
rect 577306 682638 578930 682648
rect 577306 678568 578930 678578
rect 177118 616208 180320 616562
rect 177118 616202 252734 616208
rect 253606 616202 253900 616212
rect 177118 615898 253606 616202
rect 177140 613076 253606 615898
rect 252470 613064 253606 613076
rect 253900 613064 257426 616202
rect 253606 613044 253900 613054
rect 570064 594490 570456 657162
rect 570062 594480 570460 594490
rect 121814 593602 195218 594118
rect 570062 593908 570460 593918
rect 121814 593592 259020 593602
rect 121814 593088 258596 593592
rect 121814 593086 259020 593088
rect 121814 592296 195218 593086
rect 258596 593078 259020 593086
rect 250950 592644 251150 592654
rect 571898 592644 572242 592646
rect 251150 592422 572242 592644
rect 250950 592412 251150 592422
rect 64902 591564 66344 591576
rect 252198 591564 252436 591574
rect 64902 590848 252198 591564
rect 252436 590848 252450 591564
rect 61502 536716 61792 536726
rect 32236 536484 61502 536716
rect 61502 536472 61792 536482
rect 10336 500976 12198 500986
rect 10336 499338 12198 499348
rect 64902 209704 66344 590848
rect 252198 590838 252436 590848
rect 570068 590200 570462 590206
rect 247854 590196 570462 590200
rect 247854 589926 570068 590196
rect 247858 587662 248062 589926
rect 570068 589910 570462 589920
rect 247858 587450 248062 587460
rect 224660 587298 227262 587308
rect 250604 587296 250804 587306
rect 246604 587294 250604 587296
rect 227262 587146 250604 587294
rect 224660 587136 250604 587146
rect 224662 587098 250604 587136
rect 246604 587096 250604 587098
rect 250604 587086 250804 587096
rect 251276 587296 251476 587306
rect 247246 586474 247576 586484
rect 249004 586474 249250 586482
rect 247576 586472 249250 586474
rect 247576 586274 249004 586472
rect 247246 586264 247576 586274
rect 249004 586264 249250 586274
rect 79366 585502 79672 585510
rect 250958 585502 251176 585512
rect 79366 585500 250958 585502
rect 79672 585256 250958 585500
rect 251276 585488 251476 587096
rect 251856 587286 252056 587296
rect 251856 585534 252056 587086
rect 252472 587284 252672 587294
rect 79366 585244 79672 585254
rect 250958 585246 251176 585256
rect 251280 557614 251474 585488
rect 71970 536694 72312 536704
rect 251280 536694 251476 557614
rect 72312 536484 251476 536694
rect 71970 536478 251476 536484
rect 71970 536474 72312 536478
rect 75794 500960 78128 500964
rect 251854 500960 252058 585534
rect 252472 585280 252672 587084
rect 258598 585284 259018 585294
rect 255232 585280 258598 585282
rect 252460 585098 258598 585280
rect 255232 585094 258598 585098
rect 258598 585080 259018 585090
rect 571898 555308 572242 592422
rect 571898 542534 572242 542752
rect 75782 500954 252198 500960
rect 75782 499350 75794 500954
rect 78128 499350 252198 500954
rect 75782 499312 252198 499350
rect 7640 209006 66344 209704
rect 7640 205536 8146 209006
rect 10574 205536 66344 209006
rect 7640 205064 66344 205536
rect 7640 205032 66294 205064
rect 566304 195368 567232 195378
rect 566304 182646 567232 182656
rect 572678 151048 573596 151058
rect 572678 137836 573596 137846
<< via2 >>
rect 229326 699376 230220 699750
rect 16760 696930 19950 698414
rect 10510 680624 11920 685002
rect 18390 559876 24696 563802
rect 70200 694638 71346 696412
rect 177698 695890 179686 697256
rect 570110 697722 570364 698478
rect 319098 696784 323672 697144
rect 122082 692996 123324 694248
rect 577306 678578 578930 682638
rect 571898 542752 572242 555308
rect 8146 205536 10574 209006
rect 566304 182656 567232 195368
rect 572678 137846 573596 151048
<< metal3 >>
rect 16192 698414 21160 702988
rect 16192 696930 16760 698414
rect 19950 696930 21160 698414
rect 16192 696078 21160 696930
rect 68194 696772 73202 702300
rect 68194 696766 73206 696772
rect 68204 696412 73206 696766
rect 68204 694638 70200 696412
rect 71346 694638 73206 696412
rect 68204 694296 73206 694638
rect 120194 694248 125192 702300
rect 165600 701324 170580 703066
rect 175886 701324 180874 703610
rect 165600 698698 180892 701324
rect 217294 701086 222282 703194
rect 227596 701086 232620 702386
rect 217294 699750 232620 701086
rect 217294 699376 229326 699750
rect 230220 699376 232620 699750
rect 217294 699324 232620 699376
rect 227596 699318 232620 699324
rect 318994 698830 323850 702402
rect 329290 698830 334328 702574
rect 175886 697256 180874 698698
rect 175886 695890 177698 697256
rect 179686 695890 180874 697256
rect 318994 697144 334328 698830
rect 566596 698478 571604 702996
rect 566596 697722 570110 698478
rect 570364 697722 571604 698478
rect 566596 697628 571604 697722
rect 318994 696784 319098 697144
rect 323672 696784 334328 697144
rect 318994 696682 334328 696784
rect 318994 696614 334260 696682
rect 175886 695414 180874 695890
rect 120194 692996 122082 694248
rect 123324 692996 125192 694248
rect 120194 692842 125192 692996
rect 1700 685002 12154 685242
rect 1700 680624 10510 685002
rect 11920 680624 12154 685002
rect 1700 680216 12154 680624
rect 576680 682638 583646 683014
rect 576680 678578 577306 682638
rect 578930 678578 583646 682638
rect 576680 677922 583646 678578
rect 1660 563802 25444 564242
rect 1660 559876 18390 563802
rect 24696 559876 25444 563802
rect 1660 559452 25444 559876
rect 1660 549442 5548 559452
rect 571888 555308 572252 555313
rect 571888 542752 571898 555308
rect 572242 542752 583684 555308
rect 571888 542747 572252 542752
rect 260 209688 5838 219686
rect 260 209006 11114 209688
rect 260 205536 8146 209006
rect 10574 205536 11114 209006
rect 260 204914 11114 205536
rect 1660 204888 11114 204914
rect 565826 195368 583454 196228
rect 565826 182656 566304 195368
rect 567232 182656 583454 195368
rect 565826 181378 583454 182656
rect 572370 151048 583364 151558
rect 572370 137846 572678 151048
rect 573596 137846 583364 151048
rect 572370 137130 583364 137846
use ulqc_ldo  ulqc_ldo_0
timestamp 1695692044
transform 1 0 -4393330 0 1 1242836
box 2442 -2542 5374 -645
use user_analog_proj_example  user_analog_proj_example_0
timestamp 1695692044
transform 1 0 245230 0 1 578608
box 5008 7668 7940 9565
use user_analog_project_wrapper_empty  user_analog_project_wrapper_empty_0
timestamp 1632839657
transform 1 0 0 0 1 0
box -800 -800 584800 704800
<< end >>
