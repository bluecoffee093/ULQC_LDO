magic
tech sky130A
magscale 1 2
timestamp 1699006903
<< metal2 >>
rect -2065 15292 1910 15293
rect 2502 15292 12324 15293
rect -2065 13834 12324 15292
rect -833 13833 3142 13834
rect -700 12951 280 12961
rect -700 12628 280 12638
rect 11200 12951 12180 12961
rect 11200 12628 12180 12638
rect -1909 11641 125 11959
rect -1980 9587 441 9905
rect 10250 8570 10720 8586
rect 11150 8570 11430 8580
rect 10250 8470 10260 8570
rect 10700 8478 10720 8570
rect 10700 8443 11694 8478
rect 10260 8270 10700 8280
rect 11150 8270 11430 8280
<< via2 >>
rect -700 12638 280 12951
rect 11200 12638 12180 12951
rect 10260 8280 10700 8570
<< metal3 >>
rect 470 23200 480 26999
rect 1460 23200 1470 26999
rect 10010 23200 10020 26999
rect 11000 23200 11010 26999
rect -710 12951 290 12956
rect -710 12638 -700 12951
rect 280 12638 290 12951
rect -710 12633 290 12638
rect -700 3707 280 12633
rect 480 10573 1460 23200
rect 10020 10573 11000 23200
rect 11190 12951 12190 12956
rect 11190 12638 11200 12951
rect 12180 12638 12190 12951
rect 11190 12633 12190 12638
rect 470 10273 480 10573
rect 1460 10273 1470 10573
rect 10010 10273 10020 10573
rect 11000 10273 11010 10573
rect 480 10270 1460 10273
rect 10020 10270 11000 10273
rect 10250 8570 10710 8575
rect 10250 8280 10260 8570
rect 10700 8280 10710 8570
rect 10250 8275 10710 8280
rect 11200 3708 12180 12633
rect -711 -4292 -701 3707
rect 279 -4292 289 3707
rect 11190 -4291 11200 3708
rect 12180 -4291 12190 3708
<< via3 >>
rect 480 23200 1460 26999
rect 10020 23200 11000 26999
rect 480 10273 1460 10573
rect 10020 10273 11000 10573
rect 10260 8280 10700 8570
rect -701 -4292 279 3707
rect 11200 -4291 12180 3708
<< metal4 >>
rect 470 26999 13000 27000
rect 470 23200 480 26999
rect 1460 23200 10020 26999
rect 11000 23200 13000 26999
rect 479 23199 1461 23200
rect 10019 23199 11001 23200
rect 479 10573 1461 10574
rect 479 10273 480 10573
rect 1460 10273 1461 10573
rect 479 10272 1461 10273
rect 10019 10573 11001 10574
rect 10019 10273 10020 10573
rect 11000 10273 11001 10573
rect 10019 10272 11001 10273
rect 10250 8570 10720 8586
rect 10250 8280 10260 8570
rect 10700 8478 10720 8570
rect 10700 8280 12320 8478
rect 10250 8240 12320 8280
rect 10250 7764 11710 8240
rect 10250 7600 12320 7764
rect 10250 7590 11695 7600
rect 11199 3708 12181 3709
rect -702 3707 11200 3708
rect -702 -4292 -701 3707
rect 279 -4291 11200 3707
rect 12180 -4291 12181 3708
rect 279 -4292 12181 -4291
rect -702 -4293 280 -4292
<< metal5 >>
rect 34251 27068 42251 31068
rect 42651 22784 50651 31068
use opamp  opamp_0
timestamp 1698954266
transform 1 0 4974 0 1 11572
box -4984 -11574 6608 2262
use power_transistor  power_transistor_0
timestamp 1699006509
transform 1 0 12633 0 1 -2709
box -938 -8491 38018 29797
<< labels >>
flabel metal4 3521 -3806 9138 -1800 0 FreeSans 8000 0 0 0 VSS
port 2 nsew
flabel metal5 34251 27068 42251 31068 0 FreeSans 8000 0 0 0 VIN
port 1 nsew
flabel metal5 42651 27067 50651 31068 0 FreeSans 8000 0 0 0 OUT
port 6 nsew
flabel metal2 -1980 9587 -1552 9905 0 FreeSans 3200 0 0 0 BGR_IN
port 4 nsew
flabel metal2 -1909 11641 -1481 11959 0 FreeSans 3200 0 0 0 ADJ
port 3 nsew
flabel metal2 -2065 13834 -721 15293 0 FreeSans 3200 0 0 0 EA_OUT
port 5 nsew
<< end >>
