magic
tech sky130A
magscale 1 2
timestamp 1697921354
<< nwell >>
rect -130 -127 21946 21433
<< psubdiff >>
rect -190 21459 22006 21493
rect -190 -153 -156 21459
rect 21972 -153 22006 21459
rect -190 -187 22006 -153
<< nsubdiff >>
rect -94 21363 21910 21397
rect -94 -57 -60 21363
rect 1630 21194 1708 21221
rect 1630 20791 1708 20818
rect 3458 21194 3536 21221
rect 3458 20791 3536 20818
rect 5286 21194 5364 21221
rect 5286 20791 5364 20818
rect 7114 21194 7192 21221
rect 7114 20791 7192 20818
rect 8942 21194 9020 21221
rect 8942 20791 9020 20818
rect 10770 21194 10848 21221
rect 10770 20791 10848 20818
rect 12598 21194 12676 21221
rect 12598 20791 12676 20818
rect 14426 21194 14504 21221
rect 14426 20791 14504 20818
rect 16254 21194 16332 21221
rect 16254 20791 16332 20818
rect 18082 21194 18160 21221
rect 18082 20791 18160 20818
rect 19910 21194 19988 21221
rect 19910 20791 19988 20818
rect 21738 21194 21816 21221
rect 21738 20791 21816 20818
rect 1630 20480 1708 20507
rect 1630 20077 1708 20104
rect 3458 20480 3536 20507
rect 3458 20077 3536 20104
rect 5286 20480 5364 20507
rect 5286 20077 5364 20104
rect 7114 20480 7192 20507
rect 7114 20077 7192 20104
rect 8942 20480 9020 20507
rect 8942 20077 9020 20104
rect 10770 20480 10848 20507
rect 10770 20077 10848 20104
rect 12598 20480 12676 20507
rect 12598 20077 12676 20104
rect 14426 20480 14504 20507
rect 14426 20077 14504 20104
rect 16254 20480 16332 20507
rect 16254 20077 16332 20104
rect 18082 20480 18160 20507
rect 18082 20077 18160 20104
rect 19910 20480 19988 20507
rect 19910 20077 19988 20104
rect 21738 20480 21816 20507
rect 21738 20077 21816 20104
rect 1630 19766 1708 19793
rect 1630 19363 1708 19390
rect 3458 19766 3536 19793
rect 3458 19363 3536 19390
rect 5286 19766 5364 19793
rect 5286 19363 5364 19390
rect 7114 19766 7192 19793
rect 7114 19363 7192 19390
rect 8942 19766 9020 19793
rect 8942 19363 9020 19390
rect 10770 19766 10848 19793
rect 10770 19363 10848 19390
rect 12598 19766 12676 19793
rect 12598 19363 12676 19390
rect 14426 19766 14504 19793
rect 14426 19363 14504 19390
rect 16254 19766 16332 19793
rect 16254 19363 16332 19390
rect 18082 19766 18160 19793
rect 18082 19363 18160 19390
rect 19910 19766 19988 19793
rect 19910 19363 19988 19390
rect 21738 19766 21816 19793
rect 21738 19363 21816 19390
rect 1630 19052 1708 19079
rect 1630 18649 1708 18676
rect 3458 19052 3536 19079
rect 3458 18649 3536 18676
rect 5286 19052 5364 19079
rect 5286 18649 5364 18676
rect 7114 19052 7192 19079
rect 7114 18649 7192 18676
rect 8942 19052 9020 19079
rect 8942 18649 9020 18676
rect 10770 19052 10848 19079
rect 10770 18649 10848 18676
rect 12598 19052 12676 19079
rect 12598 18649 12676 18676
rect 14426 19052 14504 19079
rect 14426 18649 14504 18676
rect 16254 19052 16332 19079
rect 16254 18649 16332 18676
rect 18082 19052 18160 19079
rect 18082 18649 18160 18676
rect 19910 19052 19988 19079
rect 19910 18649 19988 18676
rect 21738 19052 21816 19079
rect 21738 18649 21816 18676
rect 1630 18338 1708 18365
rect 1630 17935 1708 17962
rect 3458 18338 3536 18365
rect 3458 17935 3536 17962
rect 5286 18338 5364 18365
rect 5286 17935 5364 17962
rect 7114 18338 7192 18365
rect 7114 17935 7192 17962
rect 8942 18338 9020 18365
rect 8942 17935 9020 17962
rect 10770 18338 10848 18365
rect 10770 17935 10848 17962
rect 12598 18338 12676 18365
rect 12598 17935 12676 17962
rect 14426 18338 14504 18365
rect 14426 17935 14504 17962
rect 16254 18338 16332 18365
rect 16254 17935 16332 17962
rect 18082 18338 18160 18365
rect 18082 17935 18160 17962
rect 19910 18338 19988 18365
rect 19910 17935 19988 17962
rect 21738 18338 21816 18365
rect 21738 17935 21816 17962
rect 1630 17624 1708 17651
rect 1630 17221 1708 17248
rect 3458 17624 3536 17651
rect 3458 17221 3536 17248
rect 5286 17624 5364 17651
rect 5286 17221 5364 17248
rect 7114 17624 7192 17651
rect 7114 17221 7192 17248
rect 8942 17624 9020 17651
rect 8942 17221 9020 17248
rect 10770 17624 10848 17651
rect 10770 17221 10848 17248
rect 12598 17624 12676 17651
rect 12598 17221 12676 17248
rect 14426 17624 14504 17651
rect 14426 17221 14504 17248
rect 16254 17624 16332 17651
rect 16254 17221 16332 17248
rect 18082 17624 18160 17651
rect 18082 17221 18160 17248
rect 19910 17624 19988 17651
rect 19910 17221 19988 17248
rect 21738 17624 21816 17651
rect 21738 17221 21816 17248
rect 1630 16910 1708 16937
rect 1630 16507 1708 16534
rect 3458 16910 3536 16937
rect 3458 16507 3536 16534
rect 5286 16910 5364 16937
rect 5286 16507 5364 16534
rect 7114 16910 7192 16937
rect 7114 16507 7192 16534
rect 8942 16910 9020 16937
rect 8942 16507 9020 16534
rect 10770 16910 10848 16937
rect 10770 16507 10848 16534
rect 12598 16910 12676 16937
rect 12598 16507 12676 16534
rect 14426 16910 14504 16937
rect 14426 16507 14504 16534
rect 16254 16910 16332 16937
rect 16254 16507 16332 16534
rect 18082 16910 18160 16937
rect 18082 16507 18160 16534
rect 19910 16910 19988 16937
rect 19910 16507 19988 16534
rect 21738 16910 21816 16937
rect 21738 16507 21816 16534
rect 1630 16196 1708 16223
rect 1630 15793 1708 15820
rect 3458 16196 3536 16223
rect 3458 15793 3536 15820
rect 5286 16196 5364 16223
rect 5286 15793 5364 15820
rect 7114 16196 7192 16223
rect 7114 15793 7192 15820
rect 8942 16196 9020 16223
rect 8942 15793 9020 15820
rect 10770 16196 10848 16223
rect 10770 15793 10848 15820
rect 12598 16196 12676 16223
rect 12598 15793 12676 15820
rect 14426 16196 14504 16223
rect 14426 15793 14504 15820
rect 16254 16196 16332 16223
rect 16254 15793 16332 15820
rect 18082 16196 18160 16223
rect 18082 15793 18160 15820
rect 19910 16196 19988 16223
rect 19910 15793 19988 15820
rect 21738 16196 21816 16223
rect 21738 15793 21816 15820
rect 1630 15482 1708 15509
rect 1630 15079 1708 15106
rect 3458 15482 3536 15509
rect 3458 15079 3536 15106
rect 5286 15482 5364 15509
rect 5286 15079 5364 15106
rect 7114 15482 7192 15509
rect 7114 15079 7192 15106
rect 8942 15482 9020 15509
rect 8942 15079 9020 15106
rect 10770 15482 10848 15509
rect 10770 15079 10848 15106
rect 12598 15482 12676 15509
rect 12598 15079 12676 15106
rect 14426 15482 14504 15509
rect 14426 15079 14504 15106
rect 16254 15482 16332 15509
rect 16254 15079 16332 15106
rect 18082 15482 18160 15509
rect 18082 15079 18160 15106
rect 19910 15482 19988 15509
rect 19910 15079 19988 15106
rect 21738 15482 21816 15509
rect 21738 15079 21816 15106
rect 1630 14768 1708 14795
rect 1630 14365 1708 14392
rect 3458 14768 3536 14795
rect 3458 14365 3536 14392
rect 5286 14768 5364 14795
rect 5286 14365 5364 14392
rect 7114 14768 7192 14795
rect 7114 14365 7192 14392
rect 8942 14768 9020 14795
rect 8942 14365 9020 14392
rect 10770 14768 10848 14795
rect 10770 14365 10848 14392
rect 12598 14768 12676 14795
rect 12598 14365 12676 14392
rect 14426 14768 14504 14795
rect 14426 14365 14504 14392
rect 16254 14768 16332 14795
rect 16254 14365 16332 14392
rect 18082 14768 18160 14795
rect 18082 14365 18160 14392
rect 19910 14768 19988 14795
rect 19910 14365 19988 14392
rect 21738 14768 21816 14795
rect 21738 14365 21816 14392
rect 1630 14054 1708 14081
rect 1630 13651 1708 13678
rect 3458 14054 3536 14081
rect 3458 13651 3536 13678
rect 5286 14054 5364 14081
rect 5286 13651 5364 13678
rect 7114 14054 7192 14081
rect 7114 13651 7192 13678
rect 8942 14054 9020 14081
rect 8942 13651 9020 13678
rect 10770 14054 10848 14081
rect 10770 13651 10848 13678
rect 12598 14054 12676 14081
rect 12598 13651 12676 13678
rect 14426 14054 14504 14081
rect 14426 13651 14504 13678
rect 16254 14054 16332 14081
rect 16254 13651 16332 13678
rect 18082 14054 18160 14081
rect 18082 13651 18160 13678
rect 19910 14054 19988 14081
rect 19910 13651 19988 13678
rect 21738 14054 21816 14081
rect 21738 13651 21816 13678
rect 1630 13340 1708 13367
rect 1630 12937 1708 12964
rect 3458 13340 3536 13367
rect 3458 12937 3536 12964
rect 5286 13340 5364 13367
rect 5286 12937 5364 12964
rect 7114 13340 7192 13367
rect 7114 12937 7192 12964
rect 8942 13340 9020 13367
rect 8942 12937 9020 12964
rect 10770 13340 10848 13367
rect 10770 12937 10848 12964
rect 12598 13340 12676 13367
rect 12598 12937 12676 12964
rect 14426 13340 14504 13367
rect 14426 12937 14504 12964
rect 16254 13340 16332 13367
rect 16254 12937 16332 12964
rect 18082 13340 18160 13367
rect 18082 12937 18160 12964
rect 19910 13340 19988 13367
rect 19910 12937 19988 12964
rect 21738 13340 21816 13367
rect 21738 12937 21816 12964
rect 1630 12626 1708 12653
rect 1630 12223 1708 12250
rect 3458 12626 3536 12653
rect 3458 12223 3536 12250
rect 5286 12626 5364 12653
rect 5286 12223 5364 12250
rect 7114 12626 7192 12653
rect 7114 12223 7192 12250
rect 8942 12626 9020 12653
rect 8942 12223 9020 12250
rect 10770 12626 10848 12653
rect 10770 12223 10848 12250
rect 12598 12626 12676 12653
rect 12598 12223 12676 12250
rect 14426 12626 14504 12653
rect 14426 12223 14504 12250
rect 16254 12626 16332 12653
rect 16254 12223 16332 12250
rect 18082 12626 18160 12653
rect 18082 12223 18160 12250
rect 19910 12626 19988 12653
rect 19910 12223 19988 12250
rect 21738 12626 21816 12653
rect 21738 12223 21816 12250
rect 1630 11912 1708 11939
rect 1630 11509 1708 11536
rect 3458 11912 3536 11939
rect 3458 11509 3536 11536
rect 5286 11912 5364 11939
rect 5286 11509 5364 11536
rect 7114 11912 7192 11939
rect 7114 11509 7192 11536
rect 8942 11912 9020 11939
rect 8942 11509 9020 11536
rect 10770 11912 10848 11939
rect 10770 11509 10848 11536
rect 12598 11912 12676 11939
rect 12598 11509 12676 11536
rect 14426 11912 14504 11939
rect 14426 11509 14504 11536
rect 16254 11912 16332 11939
rect 16254 11509 16332 11536
rect 18082 11912 18160 11939
rect 18082 11509 18160 11536
rect 19910 11912 19988 11939
rect 19910 11509 19988 11536
rect 21738 11912 21816 11939
rect 21738 11509 21816 11536
rect 1630 11198 1708 11225
rect 1630 10795 1708 10822
rect 3458 11198 3536 11225
rect 3458 10795 3536 10822
rect 5286 11198 5364 11225
rect 5286 10795 5364 10822
rect 7114 11198 7192 11225
rect 7114 10795 7192 10822
rect 8942 11198 9020 11225
rect 8942 10795 9020 10822
rect 10770 11198 10848 11225
rect 10770 10795 10848 10822
rect 12598 11198 12676 11225
rect 12598 10795 12676 10822
rect 14426 11198 14504 11225
rect 14426 10795 14504 10822
rect 16254 11198 16332 11225
rect 16254 10795 16332 10822
rect 18082 11198 18160 11225
rect 18082 10795 18160 10822
rect 19910 11198 19988 11225
rect 19910 10795 19988 10822
rect 21738 11198 21816 11225
rect 21738 10795 21816 10822
rect 1630 10484 1708 10511
rect 1630 10081 1708 10108
rect 3458 10484 3536 10511
rect 3458 10081 3536 10108
rect 5286 10484 5364 10511
rect 5286 10081 5364 10108
rect 7114 10484 7192 10511
rect 7114 10081 7192 10108
rect 8942 10484 9020 10511
rect 8942 10081 9020 10108
rect 10770 10484 10848 10511
rect 10770 10081 10848 10108
rect 12598 10484 12676 10511
rect 12598 10081 12676 10108
rect 14426 10484 14504 10511
rect 14426 10081 14504 10108
rect 16254 10484 16332 10511
rect 16254 10081 16332 10108
rect 18082 10484 18160 10511
rect 18082 10081 18160 10108
rect 19910 10484 19988 10511
rect 19910 10081 19988 10108
rect 21738 10484 21816 10511
rect 21738 10081 21816 10108
rect 1630 9770 1708 9797
rect 1630 9367 1708 9394
rect 3458 9770 3536 9797
rect 3458 9367 3536 9394
rect 5286 9770 5364 9797
rect 5286 9367 5364 9394
rect 7114 9770 7192 9797
rect 7114 9367 7192 9394
rect 8942 9770 9020 9797
rect 8942 9367 9020 9394
rect 10770 9770 10848 9797
rect 10770 9367 10848 9394
rect 12598 9770 12676 9797
rect 12598 9367 12676 9394
rect 14426 9770 14504 9797
rect 14426 9367 14504 9394
rect 16254 9770 16332 9797
rect 16254 9367 16332 9394
rect 18082 9770 18160 9797
rect 18082 9367 18160 9394
rect 19910 9770 19988 9797
rect 19910 9367 19988 9394
rect 21738 9770 21816 9797
rect 21738 9367 21816 9394
rect 1630 9056 1708 9083
rect 1630 8653 1708 8680
rect 3458 9056 3536 9083
rect 3458 8653 3536 8680
rect 5286 9056 5364 9083
rect 5286 8653 5364 8680
rect 7114 9056 7192 9083
rect 7114 8653 7192 8680
rect 8942 9056 9020 9083
rect 8942 8653 9020 8680
rect 10770 9056 10848 9083
rect 10770 8653 10848 8680
rect 12598 9056 12676 9083
rect 12598 8653 12676 8680
rect 14426 9056 14504 9083
rect 14426 8653 14504 8680
rect 16254 9056 16332 9083
rect 16254 8653 16332 8680
rect 18082 9056 18160 9083
rect 18082 8653 18160 8680
rect 19910 9056 19988 9083
rect 19910 8653 19988 8680
rect 21738 9056 21816 9083
rect 21738 8653 21816 8680
rect 1630 8342 1708 8369
rect 1630 7939 1708 7966
rect 3458 8342 3536 8369
rect 3458 7939 3536 7966
rect 5286 8342 5364 8369
rect 5286 7939 5364 7966
rect 7114 8342 7192 8369
rect 7114 7939 7192 7966
rect 8942 8342 9020 8369
rect 8942 7939 9020 7966
rect 10770 8342 10848 8369
rect 10770 7939 10848 7966
rect 12598 8342 12676 8369
rect 12598 7939 12676 7966
rect 14426 8342 14504 8369
rect 14426 7939 14504 7966
rect 16254 8342 16332 8369
rect 16254 7939 16332 7966
rect 18082 8342 18160 8369
rect 18082 7939 18160 7966
rect 19910 8342 19988 8369
rect 19910 7939 19988 7966
rect 21738 8342 21816 8369
rect 21738 7939 21816 7966
rect 1630 7628 1708 7655
rect 1630 7225 1708 7252
rect 3458 7628 3536 7655
rect 3458 7225 3536 7252
rect 5286 7628 5364 7655
rect 5286 7225 5364 7252
rect 7114 7628 7192 7655
rect 7114 7225 7192 7252
rect 8942 7628 9020 7655
rect 8942 7225 9020 7252
rect 10770 7628 10848 7655
rect 10770 7225 10848 7252
rect 12598 7628 12676 7655
rect 12598 7225 12676 7252
rect 14426 7628 14504 7655
rect 14426 7225 14504 7252
rect 16254 7628 16332 7655
rect 16254 7225 16332 7252
rect 18082 7628 18160 7655
rect 18082 7225 18160 7252
rect 19910 7628 19988 7655
rect 19910 7225 19988 7252
rect 21738 7628 21816 7655
rect 21738 7225 21816 7252
rect 1630 6914 1708 6941
rect 1630 6511 1708 6538
rect 3458 6914 3536 6941
rect 3458 6511 3536 6538
rect 5286 6914 5364 6941
rect 5286 6511 5364 6538
rect 7114 6914 7192 6941
rect 7114 6511 7192 6538
rect 8942 6914 9020 6941
rect 8942 6511 9020 6538
rect 10770 6914 10848 6941
rect 10770 6511 10848 6538
rect 12598 6914 12676 6941
rect 12598 6511 12676 6538
rect 14426 6914 14504 6941
rect 14426 6511 14504 6538
rect 16254 6914 16332 6941
rect 16254 6511 16332 6538
rect 18082 6914 18160 6941
rect 18082 6511 18160 6538
rect 19910 6914 19988 6941
rect 19910 6511 19988 6538
rect 21738 6914 21816 6941
rect 21738 6511 21816 6538
rect 1630 6200 1708 6227
rect 1630 5797 1708 5824
rect 3458 6200 3536 6227
rect 3458 5797 3536 5824
rect 5286 6200 5364 6227
rect 5286 5797 5364 5824
rect 7114 6200 7192 6227
rect 7114 5797 7192 5824
rect 8942 6200 9020 6227
rect 8942 5797 9020 5824
rect 10770 6200 10848 6227
rect 10770 5797 10848 5824
rect 12598 6200 12676 6227
rect 12598 5797 12676 5824
rect 14426 6200 14504 6227
rect 14426 5797 14504 5824
rect 16254 6200 16332 6227
rect 16254 5797 16332 5824
rect 18082 6200 18160 6227
rect 18082 5797 18160 5824
rect 19910 6200 19988 6227
rect 19910 5797 19988 5824
rect 21738 6200 21816 6227
rect 21738 5797 21816 5824
rect 1630 5486 1708 5513
rect 1630 5083 1708 5110
rect 3458 5486 3536 5513
rect 3458 5083 3536 5110
rect 5286 5486 5364 5513
rect 5286 5083 5364 5110
rect 7114 5486 7192 5513
rect 7114 5083 7192 5110
rect 8942 5486 9020 5513
rect 8942 5083 9020 5110
rect 10770 5486 10848 5513
rect 10770 5083 10848 5110
rect 12598 5486 12676 5513
rect 12598 5083 12676 5110
rect 14426 5486 14504 5513
rect 14426 5083 14504 5110
rect 16254 5486 16332 5513
rect 16254 5083 16332 5110
rect 18082 5486 18160 5513
rect 18082 5083 18160 5110
rect 19910 5486 19988 5513
rect 19910 5083 19988 5110
rect 21738 5486 21816 5513
rect 21738 5083 21816 5110
rect 1630 4772 1708 4799
rect 1630 4369 1708 4396
rect 3458 4772 3536 4799
rect 3458 4369 3536 4396
rect 5286 4772 5364 4799
rect 5286 4369 5364 4396
rect 7114 4772 7192 4799
rect 7114 4369 7192 4396
rect 8942 4772 9020 4799
rect 8942 4369 9020 4396
rect 10770 4772 10848 4799
rect 10770 4369 10848 4396
rect 12598 4772 12676 4799
rect 12598 4369 12676 4396
rect 14426 4772 14504 4799
rect 14426 4369 14504 4396
rect 16254 4772 16332 4799
rect 16254 4369 16332 4396
rect 18082 4772 18160 4799
rect 18082 4369 18160 4396
rect 19910 4772 19988 4799
rect 19910 4369 19988 4396
rect 21738 4772 21816 4799
rect 21738 4369 21816 4396
rect 1630 4058 1708 4085
rect 1630 3655 1708 3682
rect 3458 4058 3536 4085
rect 3458 3655 3536 3682
rect 5286 4058 5364 4085
rect 5286 3655 5364 3682
rect 7114 4058 7192 4085
rect 7114 3655 7192 3682
rect 8942 4058 9020 4085
rect 8942 3655 9020 3682
rect 10770 4058 10848 4085
rect 10770 3655 10848 3682
rect 12598 4058 12676 4085
rect 12598 3655 12676 3682
rect 14426 4058 14504 4085
rect 14426 3655 14504 3682
rect 16254 4058 16332 4085
rect 16254 3655 16332 3682
rect 18082 4058 18160 4085
rect 18082 3655 18160 3682
rect 19910 4058 19988 4085
rect 19910 3655 19988 3682
rect 21738 4058 21816 4085
rect 21738 3655 21816 3682
rect 1630 3344 1708 3371
rect 1630 2941 1708 2968
rect 3458 3344 3536 3371
rect 3458 2941 3536 2968
rect 5286 3344 5364 3371
rect 5286 2941 5364 2968
rect 7114 3344 7192 3371
rect 7114 2941 7192 2968
rect 8942 3344 9020 3371
rect 8942 2941 9020 2968
rect 10770 3344 10848 3371
rect 10770 2941 10848 2968
rect 12598 3344 12676 3371
rect 12598 2941 12676 2968
rect 14426 3344 14504 3371
rect 14426 2941 14504 2968
rect 16254 3344 16332 3371
rect 16254 2941 16332 2968
rect 18082 3344 18160 3371
rect 18082 2941 18160 2968
rect 19910 3344 19988 3371
rect 19910 2941 19988 2968
rect 21738 3344 21816 3371
rect 21738 2941 21816 2968
rect 1630 2630 1708 2657
rect 1630 2227 1708 2254
rect 3458 2630 3536 2657
rect 3458 2227 3536 2254
rect 5286 2630 5364 2657
rect 5286 2227 5364 2254
rect 7114 2630 7192 2657
rect 7114 2227 7192 2254
rect 8942 2630 9020 2657
rect 8942 2227 9020 2254
rect 10770 2630 10848 2657
rect 10770 2227 10848 2254
rect 12598 2630 12676 2657
rect 12598 2227 12676 2254
rect 14426 2630 14504 2657
rect 14426 2227 14504 2254
rect 16254 2630 16332 2657
rect 16254 2227 16332 2254
rect 18082 2630 18160 2657
rect 18082 2227 18160 2254
rect 19910 2630 19988 2657
rect 19910 2227 19988 2254
rect 21738 2630 21816 2657
rect 21738 2227 21816 2254
rect 1630 1916 1708 1943
rect 1630 1513 1708 1540
rect 3458 1916 3536 1943
rect 3458 1513 3536 1540
rect 5286 1916 5364 1943
rect 5286 1513 5364 1540
rect 7114 1916 7192 1943
rect 7114 1513 7192 1540
rect 8942 1916 9020 1943
rect 8942 1513 9020 1540
rect 10770 1916 10848 1943
rect 10770 1513 10848 1540
rect 12598 1916 12676 1943
rect 12598 1513 12676 1540
rect 14426 1916 14504 1943
rect 14426 1513 14504 1540
rect 16254 1916 16332 1943
rect 16254 1513 16332 1540
rect 18082 1916 18160 1943
rect 18082 1513 18160 1540
rect 19910 1916 19988 1943
rect 19910 1513 19988 1540
rect 21738 1916 21816 1943
rect 21738 1513 21816 1540
rect 1630 1202 1708 1229
rect 1630 799 1708 826
rect 3458 1202 3536 1229
rect 3458 799 3536 826
rect 5286 1202 5364 1229
rect 5286 799 5364 826
rect 7114 1202 7192 1229
rect 7114 799 7192 826
rect 8942 1202 9020 1229
rect 8942 799 9020 826
rect 10770 1202 10848 1229
rect 10770 799 10848 826
rect 12598 1202 12676 1229
rect 12598 799 12676 826
rect 14426 1202 14504 1229
rect 14426 799 14504 826
rect 16254 1202 16332 1229
rect 16254 799 16332 826
rect 18082 1202 18160 1229
rect 18082 799 18160 826
rect 19910 1202 19988 1229
rect 19910 799 19988 826
rect 21738 1202 21816 1229
rect 21738 799 21816 826
rect 1630 488 1708 515
rect 1630 85 1708 112
rect 3458 488 3536 515
rect 3458 85 3536 112
rect 5286 488 5364 515
rect 5286 85 5364 112
rect 7114 488 7192 515
rect 7114 85 7192 112
rect 8942 488 9020 515
rect 8942 85 9020 112
rect 10770 488 10848 515
rect 10770 85 10848 112
rect 12598 488 12676 515
rect 12598 85 12676 112
rect 14426 488 14504 515
rect 14426 85 14504 112
rect 16254 488 16332 515
rect 16254 85 16332 112
rect 18082 488 18160 515
rect 18082 85 18160 112
rect 19910 488 19988 515
rect 19910 85 19988 112
rect 21738 488 21816 515
rect 21738 85 21816 112
rect 21876 -57 21910 21363
rect -94 -91 21910 -57
<< nsubdiffcont >>
rect 1630 20818 1708 21194
rect 3458 20818 3536 21194
rect 5286 20818 5364 21194
rect 7114 20818 7192 21194
rect 8942 20818 9020 21194
rect 10770 20818 10848 21194
rect 12598 20818 12676 21194
rect 14426 20818 14504 21194
rect 16254 20818 16332 21194
rect 18082 20818 18160 21194
rect 19910 20818 19988 21194
rect 21738 20818 21816 21194
rect 1630 20104 1708 20480
rect 3458 20104 3536 20480
rect 5286 20104 5364 20480
rect 7114 20104 7192 20480
rect 8942 20104 9020 20480
rect 10770 20104 10848 20480
rect 12598 20104 12676 20480
rect 14426 20104 14504 20480
rect 16254 20104 16332 20480
rect 18082 20104 18160 20480
rect 19910 20104 19988 20480
rect 21738 20104 21816 20480
rect 1630 19390 1708 19766
rect 3458 19390 3536 19766
rect 5286 19390 5364 19766
rect 7114 19390 7192 19766
rect 8942 19390 9020 19766
rect 10770 19390 10848 19766
rect 12598 19390 12676 19766
rect 14426 19390 14504 19766
rect 16254 19390 16332 19766
rect 18082 19390 18160 19766
rect 19910 19390 19988 19766
rect 21738 19390 21816 19766
rect 1630 18676 1708 19052
rect 3458 18676 3536 19052
rect 5286 18676 5364 19052
rect 7114 18676 7192 19052
rect 8942 18676 9020 19052
rect 10770 18676 10848 19052
rect 12598 18676 12676 19052
rect 14426 18676 14504 19052
rect 16254 18676 16332 19052
rect 18082 18676 18160 19052
rect 19910 18676 19988 19052
rect 21738 18676 21816 19052
rect 1630 17962 1708 18338
rect 3458 17962 3536 18338
rect 5286 17962 5364 18338
rect 7114 17962 7192 18338
rect 8942 17962 9020 18338
rect 10770 17962 10848 18338
rect 12598 17962 12676 18338
rect 14426 17962 14504 18338
rect 16254 17962 16332 18338
rect 18082 17962 18160 18338
rect 19910 17962 19988 18338
rect 21738 17962 21816 18338
rect 1630 17248 1708 17624
rect 3458 17248 3536 17624
rect 5286 17248 5364 17624
rect 7114 17248 7192 17624
rect 8942 17248 9020 17624
rect 10770 17248 10848 17624
rect 12598 17248 12676 17624
rect 14426 17248 14504 17624
rect 16254 17248 16332 17624
rect 18082 17248 18160 17624
rect 19910 17248 19988 17624
rect 21738 17248 21816 17624
rect 1630 16534 1708 16910
rect 3458 16534 3536 16910
rect 5286 16534 5364 16910
rect 7114 16534 7192 16910
rect 8942 16534 9020 16910
rect 10770 16534 10848 16910
rect 12598 16534 12676 16910
rect 14426 16534 14504 16910
rect 16254 16534 16332 16910
rect 18082 16534 18160 16910
rect 19910 16534 19988 16910
rect 21738 16534 21816 16910
rect 1630 15820 1708 16196
rect 3458 15820 3536 16196
rect 5286 15820 5364 16196
rect 7114 15820 7192 16196
rect 8942 15820 9020 16196
rect 10770 15820 10848 16196
rect 12598 15820 12676 16196
rect 14426 15820 14504 16196
rect 16254 15820 16332 16196
rect 18082 15820 18160 16196
rect 19910 15820 19988 16196
rect 21738 15820 21816 16196
rect 1630 15106 1708 15482
rect 3458 15106 3536 15482
rect 5286 15106 5364 15482
rect 7114 15106 7192 15482
rect 8942 15106 9020 15482
rect 10770 15106 10848 15482
rect 12598 15106 12676 15482
rect 14426 15106 14504 15482
rect 16254 15106 16332 15482
rect 18082 15106 18160 15482
rect 19910 15106 19988 15482
rect 21738 15106 21816 15482
rect 1630 14392 1708 14768
rect 3458 14392 3536 14768
rect 5286 14392 5364 14768
rect 7114 14392 7192 14768
rect 8942 14392 9020 14768
rect 10770 14392 10848 14768
rect 12598 14392 12676 14768
rect 14426 14392 14504 14768
rect 16254 14392 16332 14768
rect 18082 14392 18160 14768
rect 19910 14392 19988 14768
rect 21738 14392 21816 14768
rect 1630 13678 1708 14054
rect 3458 13678 3536 14054
rect 5286 13678 5364 14054
rect 7114 13678 7192 14054
rect 8942 13678 9020 14054
rect 10770 13678 10848 14054
rect 12598 13678 12676 14054
rect 14426 13678 14504 14054
rect 16254 13678 16332 14054
rect 18082 13678 18160 14054
rect 19910 13678 19988 14054
rect 21738 13678 21816 14054
rect 1630 12964 1708 13340
rect 3458 12964 3536 13340
rect 5286 12964 5364 13340
rect 7114 12964 7192 13340
rect 8942 12964 9020 13340
rect 10770 12964 10848 13340
rect 12598 12964 12676 13340
rect 14426 12964 14504 13340
rect 16254 12964 16332 13340
rect 18082 12964 18160 13340
rect 19910 12964 19988 13340
rect 21738 12964 21816 13340
rect 1630 12250 1708 12626
rect 3458 12250 3536 12626
rect 5286 12250 5364 12626
rect 7114 12250 7192 12626
rect 8942 12250 9020 12626
rect 10770 12250 10848 12626
rect 12598 12250 12676 12626
rect 14426 12250 14504 12626
rect 16254 12250 16332 12626
rect 18082 12250 18160 12626
rect 19910 12250 19988 12626
rect 21738 12250 21816 12626
rect 1630 11536 1708 11912
rect 3458 11536 3536 11912
rect 5286 11536 5364 11912
rect 7114 11536 7192 11912
rect 8942 11536 9020 11912
rect 10770 11536 10848 11912
rect 12598 11536 12676 11912
rect 14426 11536 14504 11912
rect 16254 11536 16332 11912
rect 18082 11536 18160 11912
rect 19910 11536 19988 11912
rect 21738 11536 21816 11912
rect 1630 10822 1708 11198
rect 3458 10822 3536 11198
rect 5286 10822 5364 11198
rect 7114 10822 7192 11198
rect 8942 10822 9020 11198
rect 10770 10822 10848 11198
rect 12598 10822 12676 11198
rect 14426 10822 14504 11198
rect 16254 10822 16332 11198
rect 18082 10822 18160 11198
rect 19910 10822 19988 11198
rect 21738 10822 21816 11198
rect 1630 10108 1708 10484
rect 3458 10108 3536 10484
rect 5286 10108 5364 10484
rect 7114 10108 7192 10484
rect 8942 10108 9020 10484
rect 10770 10108 10848 10484
rect 12598 10108 12676 10484
rect 14426 10108 14504 10484
rect 16254 10108 16332 10484
rect 18082 10108 18160 10484
rect 19910 10108 19988 10484
rect 21738 10108 21816 10484
rect 1630 9394 1708 9770
rect 3458 9394 3536 9770
rect 5286 9394 5364 9770
rect 7114 9394 7192 9770
rect 8942 9394 9020 9770
rect 10770 9394 10848 9770
rect 12598 9394 12676 9770
rect 14426 9394 14504 9770
rect 16254 9394 16332 9770
rect 18082 9394 18160 9770
rect 19910 9394 19988 9770
rect 21738 9394 21816 9770
rect 1630 8680 1708 9056
rect 3458 8680 3536 9056
rect 5286 8680 5364 9056
rect 7114 8680 7192 9056
rect 8942 8680 9020 9056
rect 10770 8680 10848 9056
rect 12598 8680 12676 9056
rect 14426 8680 14504 9056
rect 16254 8680 16332 9056
rect 18082 8680 18160 9056
rect 19910 8680 19988 9056
rect 21738 8680 21816 9056
rect 1630 7966 1708 8342
rect 3458 7966 3536 8342
rect 5286 7966 5364 8342
rect 7114 7966 7192 8342
rect 8942 7966 9020 8342
rect 10770 7966 10848 8342
rect 12598 7966 12676 8342
rect 14426 7966 14504 8342
rect 16254 7966 16332 8342
rect 18082 7966 18160 8342
rect 19910 7966 19988 8342
rect 21738 7966 21816 8342
rect 1630 7252 1708 7628
rect 3458 7252 3536 7628
rect 5286 7252 5364 7628
rect 7114 7252 7192 7628
rect 8942 7252 9020 7628
rect 10770 7252 10848 7628
rect 12598 7252 12676 7628
rect 14426 7252 14504 7628
rect 16254 7252 16332 7628
rect 18082 7252 18160 7628
rect 19910 7252 19988 7628
rect 21738 7252 21816 7628
rect 1630 6538 1708 6914
rect 3458 6538 3536 6914
rect 5286 6538 5364 6914
rect 7114 6538 7192 6914
rect 8942 6538 9020 6914
rect 10770 6538 10848 6914
rect 12598 6538 12676 6914
rect 14426 6538 14504 6914
rect 16254 6538 16332 6914
rect 18082 6538 18160 6914
rect 19910 6538 19988 6914
rect 21738 6538 21816 6914
rect 1630 5824 1708 6200
rect 3458 5824 3536 6200
rect 5286 5824 5364 6200
rect 7114 5824 7192 6200
rect 8942 5824 9020 6200
rect 10770 5824 10848 6200
rect 12598 5824 12676 6200
rect 14426 5824 14504 6200
rect 16254 5824 16332 6200
rect 18082 5824 18160 6200
rect 19910 5824 19988 6200
rect 21738 5824 21816 6200
rect 1630 5110 1708 5486
rect 3458 5110 3536 5486
rect 5286 5110 5364 5486
rect 7114 5110 7192 5486
rect 8942 5110 9020 5486
rect 10770 5110 10848 5486
rect 12598 5110 12676 5486
rect 14426 5110 14504 5486
rect 16254 5110 16332 5486
rect 18082 5110 18160 5486
rect 19910 5110 19988 5486
rect 21738 5110 21816 5486
rect 1630 4396 1708 4772
rect 3458 4396 3536 4772
rect 5286 4396 5364 4772
rect 7114 4396 7192 4772
rect 8942 4396 9020 4772
rect 10770 4396 10848 4772
rect 12598 4396 12676 4772
rect 14426 4396 14504 4772
rect 16254 4396 16332 4772
rect 18082 4396 18160 4772
rect 19910 4396 19988 4772
rect 21738 4396 21816 4772
rect 1630 3682 1708 4058
rect 3458 3682 3536 4058
rect 5286 3682 5364 4058
rect 7114 3682 7192 4058
rect 8942 3682 9020 4058
rect 10770 3682 10848 4058
rect 12598 3682 12676 4058
rect 14426 3682 14504 4058
rect 16254 3682 16332 4058
rect 18082 3682 18160 4058
rect 19910 3682 19988 4058
rect 21738 3682 21816 4058
rect 1630 2968 1708 3344
rect 3458 2968 3536 3344
rect 5286 2968 5364 3344
rect 7114 2968 7192 3344
rect 8942 2968 9020 3344
rect 10770 2968 10848 3344
rect 12598 2968 12676 3344
rect 14426 2968 14504 3344
rect 16254 2968 16332 3344
rect 18082 2968 18160 3344
rect 19910 2968 19988 3344
rect 21738 2968 21816 3344
rect 1630 2254 1708 2630
rect 3458 2254 3536 2630
rect 5286 2254 5364 2630
rect 7114 2254 7192 2630
rect 8942 2254 9020 2630
rect 10770 2254 10848 2630
rect 12598 2254 12676 2630
rect 14426 2254 14504 2630
rect 16254 2254 16332 2630
rect 18082 2254 18160 2630
rect 19910 2254 19988 2630
rect 21738 2254 21816 2630
rect 1630 1540 1708 1916
rect 3458 1540 3536 1916
rect 5286 1540 5364 1916
rect 7114 1540 7192 1916
rect 8942 1540 9020 1916
rect 10770 1540 10848 1916
rect 12598 1540 12676 1916
rect 14426 1540 14504 1916
rect 16254 1540 16332 1916
rect 18082 1540 18160 1916
rect 19910 1540 19988 1916
rect 21738 1540 21816 1916
rect 1630 826 1708 1202
rect 3458 826 3536 1202
rect 5286 826 5364 1202
rect 7114 826 7192 1202
rect 8942 826 9020 1202
rect 10770 826 10848 1202
rect 12598 826 12676 1202
rect 14426 826 14504 1202
rect 16254 826 16332 1202
rect 18082 826 18160 1202
rect 19910 826 19988 1202
rect 21738 826 21816 1202
rect 1630 112 1708 488
rect 3458 112 3536 488
rect 5286 112 5364 488
rect 7114 112 7192 488
rect 8942 112 9020 488
rect 10770 112 10848 488
rect 12598 112 12676 488
rect 14426 112 14504 488
rect 16254 112 16332 488
rect 18082 112 18160 488
rect 19910 112 19988 488
rect 21738 112 21816 488
<< poly >>
rect 0 21244 1490 21303
rect 1828 21244 3318 21303
rect 3656 21244 5146 21303
rect 5484 21244 6974 21303
rect 7312 21244 8802 21303
rect 9140 21244 10630 21303
rect 10968 21244 12458 21303
rect 12796 21244 14286 21303
rect 14624 21244 16114 21303
rect 16452 21244 17942 21303
rect 18280 21244 19770 21303
rect 20108 21244 21598 21303
rect 98 21232 128 21244
rect 290 21232 320 21244
rect 482 21232 512 21244
rect 674 21232 704 21244
rect 866 21232 896 21244
rect 1058 21232 1088 21244
rect 1250 21232 1280 21244
rect 1442 21232 1472 21244
rect 1926 21232 1956 21244
rect 2118 21232 2148 21244
rect 2310 21232 2340 21244
rect 2502 21232 2532 21244
rect 2694 21232 2724 21244
rect 2886 21232 2916 21244
rect 3078 21232 3108 21244
rect 3270 21232 3300 21244
rect 3754 21232 3784 21244
rect 3946 21232 3976 21244
rect 4138 21232 4168 21244
rect 4330 21232 4360 21244
rect 4522 21232 4552 21244
rect 4714 21232 4744 21244
rect 4906 21232 4936 21244
rect 5098 21232 5128 21244
rect 5582 21232 5612 21244
rect 5774 21232 5804 21244
rect 5966 21232 5996 21244
rect 6158 21232 6188 21244
rect 6350 21232 6380 21244
rect 6542 21232 6572 21244
rect 6734 21232 6764 21244
rect 6926 21232 6956 21244
rect 7410 21232 7440 21244
rect 7602 21232 7632 21244
rect 7794 21232 7824 21244
rect 7986 21232 8016 21244
rect 8178 21232 8208 21244
rect 8370 21232 8400 21244
rect 8562 21232 8592 21244
rect 8754 21232 8784 21244
rect 9238 21232 9268 21244
rect 9430 21232 9460 21244
rect 9622 21232 9652 21244
rect 9814 21232 9844 21244
rect 10006 21232 10036 21244
rect 10198 21232 10228 21244
rect 10390 21232 10420 21244
rect 10582 21232 10612 21244
rect 11066 21232 11096 21244
rect 11258 21232 11288 21244
rect 11450 21232 11480 21244
rect 11642 21232 11672 21244
rect 11834 21232 11864 21244
rect 12026 21232 12056 21244
rect 12218 21232 12248 21244
rect 12410 21232 12440 21244
rect 12894 21232 12924 21244
rect 13086 21232 13116 21244
rect 13278 21232 13308 21244
rect 13470 21232 13500 21244
rect 13662 21232 13692 21244
rect 13854 21232 13884 21244
rect 14046 21232 14076 21244
rect 14238 21232 14268 21244
rect 14722 21232 14752 21244
rect 14914 21232 14944 21244
rect 15106 21232 15136 21244
rect 15298 21232 15328 21244
rect 15490 21232 15520 21244
rect 15682 21232 15712 21244
rect 15874 21232 15904 21244
rect 16066 21232 16096 21244
rect 16550 21232 16580 21244
rect 16742 21232 16772 21244
rect 16934 21232 16964 21244
rect 17126 21232 17156 21244
rect 17318 21232 17348 21244
rect 17510 21232 17540 21244
rect 17702 21232 17732 21244
rect 17894 21232 17924 21244
rect 18378 21232 18408 21244
rect 18570 21232 18600 21244
rect 18762 21232 18792 21244
rect 18954 21232 18984 21244
rect 19146 21232 19176 21244
rect 19338 21232 19368 21244
rect 19530 21232 19560 21244
rect 19722 21232 19752 21244
rect 20206 21232 20236 21244
rect 20398 21232 20428 21244
rect 20590 21232 20620 21244
rect 20782 21232 20812 21244
rect 20974 21232 21004 21244
rect 21166 21232 21196 21244
rect 21358 21232 21388 21244
rect 21550 21232 21580 21244
rect 194 20768 224 20780
rect 386 20768 416 20780
rect 578 20768 608 20780
rect 770 20768 800 20780
rect 962 20768 992 20780
rect 1154 20768 1184 20780
rect 1346 20768 1376 20780
rect 2022 20768 2052 20780
rect 2214 20768 2244 20780
rect 2406 20768 2436 20780
rect 2598 20768 2628 20780
rect 2790 20768 2820 20780
rect 2982 20768 3012 20780
rect 3174 20768 3204 20780
rect 3850 20768 3880 20780
rect 4042 20768 4072 20780
rect 4234 20768 4264 20780
rect 4426 20768 4456 20780
rect 4618 20768 4648 20780
rect 4810 20768 4840 20780
rect 5002 20768 5032 20780
rect 5678 20768 5708 20780
rect 5870 20768 5900 20780
rect 6062 20768 6092 20780
rect 6254 20768 6284 20780
rect 6446 20768 6476 20780
rect 6638 20768 6668 20780
rect 6830 20768 6860 20780
rect 7506 20768 7536 20780
rect 7698 20768 7728 20780
rect 7890 20768 7920 20780
rect 8082 20768 8112 20780
rect 8274 20768 8304 20780
rect 8466 20768 8496 20780
rect 8658 20768 8688 20780
rect 9334 20768 9364 20780
rect 9526 20768 9556 20780
rect 9718 20768 9748 20780
rect 9910 20768 9940 20780
rect 10102 20768 10132 20780
rect 10294 20768 10324 20780
rect 10486 20768 10516 20780
rect 11162 20768 11192 20780
rect 11354 20768 11384 20780
rect 11546 20768 11576 20780
rect 11738 20768 11768 20780
rect 11930 20768 11960 20780
rect 12122 20768 12152 20780
rect 12314 20768 12344 20780
rect 12990 20768 13020 20780
rect 13182 20768 13212 20780
rect 13374 20768 13404 20780
rect 13566 20768 13596 20780
rect 13758 20768 13788 20780
rect 13950 20768 13980 20780
rect 14142 20768 14172 20780
rect 14818 20768 14848 20780
rect 15010 20768 15040 20780
rect 15202 20768 15232 20780
rect 15394 20768 15424 20780
rect 15586 20768 15616 20780
rect 15778 20768 15808 20780
rect 15970 20768 16000 20780
rect 16646 20768 16676 20780
rect 16838 20768 16868 20780
rect 17030 20768 17060 20780
rect 17222 20768 17252 20780
rect 17414 20768 17444 20780
rect 17606 20768 17636 20780
rect 17798 20768 17828 20780
rect 18474 20768 18504 20780
rect 18666 20768 18696 20780
rect 18858 20768 18888 20780
rect 19050 20768 19080 20780
rect 19242 20768 19272 20780
rect 19434 20768 19464 20780
rect 19626 20768 19656 20780
rect 20302 20768 20332 20780
rect 20494 20768 20524 20780
rect 20686 20768 20716 20780
rect 20878 20768 20908 20780
rect 21070 20768 21100 20780
rect 21262 20768 21292 20780
rect 21454 20768 21484 20780
rect 0 20709 1490 20768
rect 1828 20709 3318 20768
rect 3656 20709 5146 20768
rect 5484 20709 6974 20768
rect 7312 20709 8802 20768
rect 9140 20709 10630 20768
rect 10968 20709 12458 20768
rect 12796 20709 14286 20768
rect 14624 20709 16114 20768
rect 16452 20709 17942 20768
rect 18280 20709 19770 20768
rect 20108 20709 21598 20768
rect 0 20530 1490 20589
rect 1828 20530 3318 20589
rect 3656 20530 5146 20589
rect 5484 20530 6974 20589
rect 7312 20530 8802 20589
rect 9140 20530 10630 20589
rect 10968 20530 12458 20589
rect 12796 20530 14286 20589
rect 14624 20530 16114 20589
rect 16452 20530 17942 20589
rect 18280 20530 19770 20589
rect 20108 20530 21598 20589
rect 98 20518 128 20530
rect 290 20518 320 20530
rect 482 20518 512 20530
rect 674 20518 704 20530
rect 866 20518 896 20530
rect 1058 20518 1088 20530
rect 1250 20518 1280 20530
rect 1442 20518 1472 20530
rect 1926 20518 1956 20530
rect 2118 20518 2148 20530
rect 2310 20518 2340 20530
rect 2502 20518 2532 20530
rect 2694 20518 2724 20530
rect 2886 20518 2916 20530
rect 3078 20518 3108 20530
rect 3270 20518 3300 20530
rect 3754 20518 3784 20530
rect 3946 20518 3976 20530
rect 4138 20518 4168 20530
rect 4330 20518 4360 20530
rect 4522 20518 4552 20530
rect 4714 20518 4744 20530
rect 4906 20518 4936 20530
rect 5098 20518 5128 20530
rect 5582 20518 5612 20530
rect 5774 20518 5804 20530
rect 5966 20518 5996 20530
rect 6158 20518 6188 20530
rect 6350 20518 6380 20530
rect 6542 20518 6572 20530
rect 6734 20518 6764 20530
rect 6926 20518 6956 20530
rect 7410 20518 7440 20530
rect 7602 20518 7632 20530
rect 7794 20518 7824 20530
rect 7986 20518 8016 20530
rect 8178 20518 8208 20530
rect 8370 20518 8400 20530
rect 8562 20518 8592 20530
rect 8754 20518 8784 20530
rect 9238 20518 9268 20530
rect 9430 20518 9460 20530
rect 9622 20518 9652 20530
rect 9814 20518 9844 20530
rect 10006 20518 10036 20530
rect 10198 20518 10228 20530
rect 10390 20518 10420 20530
rect 10582 20518 10612 20530
rect 11066 20518 11096 20530
rect 11258 20518 11288 20530
rect 11450 20518 11480 20530
rect 11642 20518 11672 20530
rect 11834 20518 11864 20530
rect 12026 20518 12056 20530
rect 12218 20518 12248 20530
rect 12410 20518 12440 20530
rect 12894 20518 12924 20530
rect 13086 20518 13116 20530
rect 13278 20518 13308 20530
rect 13470 20518 13500 20530
rect 13662 20518 13692 20530
rect 13854 20518 13884 20530
rect 14046 20518 14076 20530
rect 14238 20518 14268 20530
rect 14722 20518 14752 20530
rect 14914 20518 14944 20530
rect 15106 20518 15136 20530
rect 15298 20518 15328 20530
rect 15490 20518 15520 20530
rect 15682 20518 15712 20530
rect 15874 20518 15904 20530
rect 16066 20518 16096 20530
rect 16550 20518 16580 20530
rect 16742 20518 16772 20530
rect 16934 20518 16964 20530
rect 17126 20518 17156 20530
rect 17318 20518 17348 20530
rect 17510 20518 17540 20530
rect 17702 20518 17732 20530
rect 17894 20518 17924 20530
rect 18378 20518 18408 20530
rect 18570 20518 18600 20530
rect 18762 20518 18792 20530
rect 18954 20518 18984 20530
rect 19146 20518 19176 20530
rect 19338 20518 19368 20530
rect 19530 20518 19560 20530
rect 19722 20518 19752 20530
rect 20206 20518 20236 20530
rect 20398 20518 20428 20530
rect 20590 20518 20620 20530
rect 20782 20518 20812 20530
rect 20974 20518 21004 20530
rect 21166 20518 21196 20530
rect 21358 20518 21388 20530
rect 21550 20518 21580 20530
rect 194 20054 224 20066
rect 386 20054 416 20066
rect 578 20054 608 20066
rect 770 20054 800 20066
rect 962 20054 992 20066
rect 1154 20054 1184 20066
rect 1346 20054 1376 20066
rect 2022 20054 2052 20066
rect 2214 20054 2244 20066
rect 2406 20054 2436 20066
rect 2598 20054 2628 20066
rect 2790 20054 2820 20066
rect 2982 20054 3012 20066
rect 3174 20054 3204 20066
rect 3850 20054 3880 20066
rect 4042 20054 4072 20066
rect 4234 20054 4264 20066
rect 4426 20054 4456 20066
rect 4618 20054 4648 20066
rect 4810 20054 4840 20066
rect 5002 20054 5032 20066
rect 5678 20054 5708 20066
rect 5870 20054 5900 20066
rect 6062 20054 6092 20066
rect 6254 20054 6284 20066
rect 6446 20054 6476 20066
rect 6638 20054 6668 20066
rect 6830 20054 6860 20066
rect 7506 20054 7536 20066
rect 7698 20054 7728 20066
rect 7890 20054 7920 20066
rect 8082 20054 8112 20066
rect 8274 20054 8304 20066
rect 8466 20054 8496 20066
rect 8658 20054 8688 20066
rect 9334 20054 9364 20066
rect 9526 20054 9556 20066
rect 9718 20054 9748 20066
rect 9910 20054 9940 20066
rect 10102 20054 10132 20066
rect 10294 20054 10324 20066
rect 10486 20054 10516 20066
rect 11162 20054 11192 20066
rect 11354 20054 11384 20066
rect 11546 20054 11576 20066
rect 11738 20054 11768 20066
rect 11930 20054 11960 20066
rect 12122 20054 12152 20066
rect 12314 20054 12344 20066
rect 12990 20054 13020 20066
rect 13182 20054 13212 20066
rect 13374 20054 13404 20066
rect 13566 20054 13596 20066
rect 13758 20054 13788 20066
rect 13950 20054 13980 20066
rect 14142 20054 14172 20066
rect 14818 20054 14848 20066
rect 15010 20054 15040 20066
rect 15202 20054 15232 20066
rect 15394 20054 15424 20066
rect 15586 20054 15616 20066
rect 15778 20054 15808 20066
rect 15970 20054 16000 20066
rect 16646 20054 16676 20066
rect 16838 20054 16868 20066
rect 17030 20054 17060 20066
rect 17222 20054 17252 20066
rect 17414 20054 17444 20066
rect 17606 20054 17636 20066
rect 17798 20054 17828 20066
rect 18474 20054 18504 20066
rect 18666 20054 18696 20066
rect 18858 20054 18888 20066
rect 19050 20054 19080 20066
rect 19242 20054 19272 20066
rect 19434 20054 19464 20066
rect 19626 20054 19656 20066
rect 20302 20054 20332 20066
rect 20494 20054 20524 20066
rect 20686 20054 20716 20066
rect 20878 20054 20908 20066
rect 21070 20054 21100 20066
rect 21262 20054 21292 20066
rect 21454 20054 21484 20066
rect 0 19995 1490 20054
rect 1828 19995 3318 20054
rect 3656 19995 5146 20054
rect 5484 19995 6974 20054
rect 7312 19995 8802 20054
rect 9140 19995 10630 20054
rect 10968 19995 12458 20054
rect 12796 19995 14286 20054
rect 14624 19995 16114 20054
rect 16452 19995 17942 20054
rect 18280 19995 19770 20054
rect 20108 19995 21598 20054
rect 0 19816 1490 19875
rect 1828 19816 3318 19875
rect 3656 19816 5146 19875
rect 5484 19816 6974 19875
rect 7312 19816 8802 19875
rect 9140 19816 10630 19875
rect 10968 19816 12458 19875
rect 12796 19816 14286 19875
rect 14624 19816 16114 19875
rect 16452 19816 17942 19875
rect 18280 19816 19770 19875
rect 20108 19816 21598 19875
rect 98 19804 128 19816
rect 290 19804 320 19816
rect 482 19804 512 19816
rect 674 19804 704 19816
rect 866 19804 896 19816
rect 1058 19804 1088 19816
rect 1250 19804 1280 19816
rect 1442 19804 1472 19816
rect 1926 19804 1956 19816
rect 2118 19804 2148 19816
rect 2310 19804 2340 19816
rect 2502 19804 2532 19816
rect 2694 19804 2724 19816
rect 2886 19804 2916 19816
rect 3078 19804 3108 19816
rect 3270 19804 3300 19816
rect 3754 19804 3784 19816
rect 3946 19804 3976 19816
rect 4138 19804 4168 19816
rect 4330 19804 4360 19816
rect 4522 19804 4552 19816
rect 4714 19804 4744 19816
rect 4906 19804 4936 19816
rect 5098 19804 5128 19816
rect 5582 19804 5612 19816
rect 5774 19804 5804 19816
rect 5966 19804 5996 19816
rect 6158 19804 6188 19816
rect 6350 19804 6380 19816
rect 6542 19804 6572 19816
rect 6734 19804 6764 19816
rect 6926 19804 6956 19816
rect 7410 19804 7440 19816
rect 7602 19804 7632 19816
rect 7794 19804 7824 19816
rect 7986 19804 8016 19816
rect 8178 19804 8208 19816
rect 8370 19804 8400 19816
rect 8562 19804 8592 19816
rect 8754 19804 8784 19816
rect 9238 19804 9268 19816
rect 9430 19804 9460 19816
rect 9622 19804 9652 19816
rect 9814 19804 9844 19816
rect 10006 19804 10036 19816
rect 10198 19804 10228 19816
rect 10390 19804 10420 19816
rect 10582 19804 10612 19816
rect 11066 19804 11096 19816
rect 11258 19804 11288 19816
rect 11450 19804 11480 19816
rect 11642 19804 11672 19816
rect 11834 19804 11864 19816
rect 12026 19804 12056 19816
rect 12218 19804 12248 19816
rect 12410 19804 12440 19816
rect 12894 19804 12924 19816
rect 13086 19804 13116 19816
rect 13278 19804 13308 19816
rect 13470 19804 13500 19816
rect 13662 19804 13692 19816
rect 13854 19804 13884 19816
rect 14046 19804 14076 19816
rect 14238 19804 14268 19816
rect 14722 19804 14752 19816
rect 14914 19804 14944 19816
rect 15106 19804 15136 19816
rect 15298 19804 15328 19816
rect 15490 19804 15520 19816
rect 15682 19804 15712 19816
rect 15874 19804 15904 19816
rect 16066 19804 16096 19816
rect 16550 19804 16580 19816
rect 16742 19804 16772 19816
rect 16934 19804 16964 19816
rect 17126 19804 17156 19816
rect 17318 19804 17348 19816
rect 17510 19804 17540 19816
rect 17702 19804 17732 19816
rect 17894 19804 17924 19816
rect 18378 19804 18408 19816
rect 18570 19804 18600 19816
rect 18762 19804 18792 19816
rect 18954 19804 18984 19816
rect 19146 19804 19176 19816
rect 19338 19804 19368 19816
rect 19530 19804 19560 19816
rect 19722 19804 19752 19816
rect 20206 19804 20236 19816
rect 20398 19804 20428 19816
rect 20590 19804 20620 19816
rect 20782 19804 20812 19816
rect 20974 19804 21004 19816
rect 21166 19804 21196 19816
rect 21358 19804 21388 19816
rect 21550 19804 21580 19816
rect 194 19340 224 19352
rect 386 19340 416 19352
rect 578 19340 608 19352
rect 770 19340 800 19352
rect 962 19340 992 19352
rect 1154 19340 1184 19352
rect 1346 19340 1376 19352
rect 2022 19340 2052 19352
rect 2214 19340 2244 19352
rect 2406 19340 2436 19352
rect 2598 19340 2628 19352
rect 2790 19340 2820 19352
rect 2982 19340 3012 19352
rect 3174 19340 3204 19352
rect 3850 19340 3880 19352
rect 4042 19340 4072 19352
rect 4234 19340 4264 19352
rect 4426 19340 4456 19352
rect 4618 19340 4648 19352
rect 4810 19340 4840 19352
rect 5002 19340 5032 19352
rect 5678 19340 5708 19352
rect 5870 19340 5900 19352
rect 6062 19340 6092 19352
rect 6254 19340 6284 19352
rect 6446 19340 6476 19352
rect 6638 19340 6668 19352
rect 6830 19340 6860 19352
rect 7506 19340 7536 19352
rect 7698 19340 7728 19352
rect 7890 19340 7920 19352
rect 8082 19340 8112 19352
rect 8274 19340 8304 19352
rect 8466 19340 8496 19352
rect 8658 19340 8688 19352
rect 9334 19340 9364 19352
rect 9526 19340 9556 19352
rect 9718 19340 9748 19352
rect 9910 19340 9940 19352
rect 10102 19340 10132 19352
rect 10294 19340 10324 19352
rect 10486 19340 10516 19352
rect 11162 19340 11192 19352
rect 11354 19340 11384 19352
rect 11546 19340 11576 19352
rect 11738 19340 11768 19352
rect 11930 19340 11960 19352
rect 12122 19340 12152 19352
rect 12314 19340 12344 19352
rect 12990 19340 13020 19352
rect 13182 19340 13212 19352
rect 13374 19340 13404 19352
rect 13566 19340 13596 19352
rect 13758 19340 13788 19352
rect 13950 19340 13980 19352
rect 14142 19340 14172 19352
rect 14818 19340 14848 19352
rect 15010 19340 15040 19352
rect 15202 19340 15232 19352
rect 15394 19340 15424 19352
rect 15586 19340 15616 19352
rect 15778 19340 15808 19352
rect 15970 19340 16000 19352
rect 16646 19340 16676 19352
rect 16838 19340 16868 19352
rect 17030 19340 17060 19352
rect 17222 19340 17252 19352
rect 17414 19340 17444 19352
rect 17606 19340 17636 19352
rect 17798 19340 17828 19352
rect 18474 19340 18504 19352
rect 18666 19340 18696 19352
rect 18858 19340 18888 19352
rect 19050 19340 19080 19352
rect 19242 19340 19272 19352
rect 19434 19340 19464 19352
rect 19626 19340 19656 19352
rect 20302 19340 20332 19352
rect 20494 19340 20524 19352
rect 20686 19340 20716 19352
rect 20878 19340 20908 19352
rect 21070 19340 21100 19352
rect 21262 19340 21292 19352
rect 21454 19340 21484 19352
rect 0 19281 1490 19340
rect 1828 19281 3318 19340
rect 3656 19281 5146 19340
rect 5484 19281 6974 19340
rect 7312 19281 8802 19340
rect 9140 19281 10630 19340
rect 10968 19281 12458 19340
rect 12796 19281 14286 19340
rect 14624 19281 16114 19340
rect 16452 19281 17942 19340
rect 18280 19281 19770 19340
rect 20108 19281 21598 19340
rect 0 19102 1490 19161
rect 1828 19102 3318 19161
rect 3656 19102 5146 19161
rect 5484 19102 6974 19161
rect 7312 19102 8802 19161
rect 9140 19102 10630 19161
rect 10968 19102 12458 19161
rect 12796 19102 14286 19161
rect 14624 19102 16114 19161
rect 16452 19102 17942 19161
rect 18280 19102 19770 19161
rect 20108 19102 21598 19161
rect 98 19090 128 19102
rect 290 19090 320 19102
rect 482 19090 512 19102
rect 674 19090 704 19102
rect 866 19090 896 19102
rect 1058 19090 1088 19102
rect 1250 19090 1280 19102
rect 1442 19090 1472 19102
rect 1926 19090 1956 19102
rect 2118 19090 2148 19102
rect 2310 19090 2340 19102
rect 2502 19090 2532 19102
rect 2694 19090 2724 19102
rect 2886 19090 2916 19102
rect 3078 19090 3108 19102
rect 3270 19090 3300 19102
rect 3754 19090 3784 19102
rect 3946 19090 3976 19102
rect 4138 19090 4168 19102
rect 4330 19090 4360 19102
rect 4522 19090 4552 19102
rect 4714 19090 4744 19102
rect 4906 19090 4936 19102
rect 5098 19090 5128 19102
rect 5582 19090 5612 19102
rect 5774 19090 5804 19102
rect 5966 19090 5996 19102
rect 6158 19090 6188 19102
rect 6350 19090 6380 19102
rect 6542 19090 6572 19102
rect 6734 19090 6764 19102
rect 6926 19090 6956 19102
rect 7410 19090 7440 19102
rect 7602 19090 7632 19102
rect 7794 19090 7824 19102
rect 7986 19090 8016 19102
rect 8178 19090 8208 19102
rect 8370 19090 8400 19102
rect 8562 19090 8592 19102
rect 8754 19090 8784 19102
rect 9238 19090 9268 19102
rect 9430 19090 9460 19102
rect 9622 19090 9652 19102
rect 9814 19090 9844 19102
rect 10006 19090 10036 19102
rect 10198 19090 10228 19102
rect 10390 19090 10420 19102
rect 10582 19090 10612 19102
rect 11066 19090 11096 19102
rect 11258 19090 11288 19102
rect 11450 19090 11480 19102
rect 11642 19090 11672 19102
rect 11834 19090 11864 19102
rect 12026 19090 12056 19102
rect 12218 19090 12248 19102
rect 12410 19090 12440 19102
rect 12894 19090 12924 19102
rect 13086 19090 13116 19102
rect 13278 19090 13308 19102
rect 13470 19090 13500 19102
rect 13662 19090 13692 19102
rect 13854 19090 13884 19102
rect 14046 19090 14076 19102
rect 14238 19090 14268 19102
rect 14722 19090 14752 19102
rect 14914 19090 14944 19102
rect 15106 19090 15136 19102
rect 15298 19090 15328 19102
rect 15490 19090 15520 19102
rect 15682 19090 15712 19102
rect 15874 19090 15904 19102
rect 16066 19090 16096 19102
rect 16550 19090 16580 19102
rect 16742 19090 16772 19102
rect 16934 19090 16964 19102
rect 17126 19090 17156 19102
rect 17318 19090 17348 19102
rect 17510 19090 17540 19102
rect 17702 19090 17732 19102
rect 17894 19090 17924 19102
rect 18378 19090 18408 19102
rect 18570 19090 18600 19102
rect 18762 19090 18792 19102
rect 18954 19090 18984 19102
rect 19146 19090 19176 19102
rect 19338 19090 19368 19102
rect 19530 19090 19560 19102
rect 19722 19090 19752 19102
rect 20206 19090 20236 19102
rect 20398 19090 20428 19102
rect 20590 19090 20620 19102
rect 20782 19090 20812 19102
rect 20974 19090 21004 19102
rect 21166 19090 21196 19102
rect 21358 19090 21388 19102
rect 21550 19090 21580 19102
rect 194 18626 224 18638
rect 386 18626 416 18638
rect 578 18626 608 18638
rect 770 18626 800 18638
rect 962 18626 992 18638
rect 1154 18626 1184 18638
rect 1346 18626 1376 18638
rect 2022 18626 2052 18638
rect 2214 18626 2244 18638
rect 2406 18626 2436 18638
rect 2598 18626 2628 18638
rect 2790 18626 2820 18638
rect 2982 18626 3012 18638
rect 3174 18626 3204 18638
rect 3850 18626 3880 18638
rect 4042 18626 4072 18638
rect 4234 18626 4264 18638
rect 4426 18626 4456 18638
rect 4618 18626 4648 18638
rect 4810 18626 4840 18638
rect 5002 18626 5032 18638
rect 5678 18626 5708 18638
rect 5870 18626 5900 18638
rect 6062 18626 6092 18638
rect 6254 18626 6284 18638
rect 6446 18626 6476 18638
rect 6638 18626 6668 18638
rect 6830 18626 6860 18638
rect 7506 18626 7536 18638
rect 7698 18626 7728 18638
rect 7890 18626 7920 18638
rect 8082 18626 8112 18638
rect 8274 18626 8304 18638
rect 8466 18626 8496 18638
rect 8658 18626 8688 18638
rect 9334 18626 9364 18638
rect 9526 18626 9556 18638
rect 9718 18626 9748 18638
rect 9910 18626 9940 18638
rect 10102 18626 10132 18638
rect 10294 18626 10324 18638
rect 10486 18626 10516 18638
rect 11162 18626 11192 18638
rect 11354 18626 11384 18638
rect 11546 18626 11576 18638
rect 11738 18626 11768 18638
rect 11930 18626 11960 18638
rect 12122 18626 12152 18638
rect 12314 18626 12344 18638
rect 12990 18626 13020 18638
rect 13182 18626 13212 18638
rect 13374 18626 13404 18638
rect 13566 18626 13596 18638
rect 13758 18626 13788 18638
rect 13950 18626 13980 18638
rect 14142 18626 14172 18638
rect 14818 18626 14848 18638
rect 15010 18626 15040 18638
rect 15202 18626 15232 18638
rect 15394 18626 15424 18638
rect 15586 18626 15616 18638
rect 15778 18626 15808 18638
rect 15970 18626 16000 18638
rect 16646 18626 16676 18638
rect 16838 18626 16868 18638
rect 17030 18626 17060 18638
rect 17222 18626 17252 18638
rect 17414 18626 17444 18638
rect 17606 18626 17636 18638
rect 17798 18626 17828 18638
rect 18474 18626 18504 18638
rect 18666 18626 18696 18638
rect 18858 18626 18888 18638
rect 19050 18626 19080 18638
rect 19242 18626 19272 18638
rect 19434 18626 19464 18638
rect 19626 18626 19656 18638
rect 20302 18626 20332 18638
rect 20494 18626 20524 18638
rect 20686 18626 20716 18638
rect 20878 18626 20908 18638
rect 21070 18626 21100 18638
rect 21262 18626 21292 18638
rect 21454 18626 21484 18638
rect 0 18567 1490 18626
rect 1828 18567 3318 18626
rect 3656 18567 5146 18626
rect 5484 18567 6974 18626
rect 7312 18567 8802 18626
rect 9140 18567 10630 18626
rect 10968 18567 12458 18626
rect 12796 18567 14286 18626
rect 14624 18567 16114 18626
rect 16452 18567 17942 18626
rect 18280 18567 19770 18626
rect 20108 18567 21598 18626
rect 0 18388 1490 18447
rect 1828 18388 3318 18447
rect 3656 18388 5146 18447
rect 5484 18388 6974 18447
rect 7312 18388 8802 18447
rect 9140 18388 10630 18447
rect 10968 18388 12458 18447
rect 12796 18388 14286 18447
rect 14624 18388 16114 18447
rect 16452 18388 17942 18447
rect 18280 18388 19770 18447
rect 20108 18388 21598 18447
rect 98 18376 128 18388
rect 290 18376 320 18388
rect 482 18376 512 18388
rect 674 18376 704 18388
rect 866 18376 896 18388
rect 1058 18376 1088 18388
rect 1250 18376 1280 18388
rect 1442 18376 1472 18388
rect 1926 18376 1956 18388
rect 2118 18376 2148 18388
rect 2310 18376 2340 18388
rect 2502 18376 2532 18388
rect 2694 18376 2724 18388
rect 2886 18376 2916 18388
rect 3078 18376 3108 18388
rect 3270 18376 3300 18388
rect 3754 18376 3784 18388
rect 3946 18376 3976 18388
rect 4138 18376 4168 18388
rect 4330 18376 4360 18388
rect 4522 18376 4552 18388
rect 4714 18376 4744 18388
rect 4906 18376 4936 18388
rect 5098 18376 5128 18388
rect 5582 18376 5612 18388
rect 5774 18376 5804 18388
rect 5966 18376 5996 18388
rect 6158 18376 6188 18388
rect 6350 18376 6380 18388
rect 6542 18376 6572 18388
rect 6734 18376 6764 18388
rect 6926 18376 6956 18388
rect 7410 18376 7440 18388
rect 7602 18376 7632 18388
rect 7794 18376 7824 18388
rect 7986 18376 8016 18388
rect 8178 18376 8208 18388
rect 8370 18376 8400 18388
rect 8562 18376 8592 18388
rect 8754 18376 8784 18388
rect 9238 18376 9268 18388
rect 9430 18376 9460 18388
rect 9622 18376 9652 18388
rect 9814 18376 9844 18388
rect 10006 18376 10036 18388
rect 10198 18376 10228 18388
rect 10390 18376 10420 18388
rect 10582 18376 10612 18388
rect 11066 18376 11096 18388
rect 11258 18376 11288 18388
rect 11450 18376 11480 18388
rect 11642 18376 11672 18388
rect 11834 18376 11864 18388
rect 12026 18376 12056 18388
rect 12218 18376 12248 18388
rect 12410 18376 12440 18388
rect 12894 18376 12924 18388
rect 13086 18376 13116 18388
rect 13278 18376 13308 18388
rect 13470 18376 13500 18388
rect 13662 18376 13692 18388
rect 13854 18376 13884 18388
rect 14046 18376 14076 18388
rect 14238 18376 14268 18388
rect 14722 18376 14752 18388
rect 14914 18376 14944 18388
rect 15106 18376 15136 18388
rect 15298 18376 15328 18388
rect 15490 18376 15520 18388
rect 15682 18376 15712 18388
rect 15874 18376 15904 18388
rect 16066 18376 16096 18388
rect 16550 18376 16580 18388
rect 16742 18376 16772 18388
rect 16934 18376 16964 18388
rect 17126 18376 17156 18388
rect 17318 18376 17348 18388
rect 17510 18376 17540 18388
rect 17702 18376 17732 18388
rect 17894 18376 17924 18388
rect 18378 18376 18408 18388
rect 18570 18376 18600 18388
rect 18762 18376 18792 18388
rect 18954 18376 18984 18388
rect 19146 18376 19176 18388
rect 19338 18376 19368 18388
rect 19530 18376 19560 18388
rect 19722 18376 19752 18388
rect 20206 18376 20236 18388
rect 20398 18376 20428 18388
rect 20590 18376 20620 18388
rect 20782 18376 20812 18388
rect 20974 18376 21004 18388
rect 21166 18376 21196 18388
rect 21358 18376 21388 18388
rect 21550 18376 21580 18388
rect 194 17912 224 17924
rect 386 17912 416 17924
rect 578 17912 608 17924
rect 770 17912 800 17924
rect 962 17912 992 17924
rect 1154 17912 1184 17924
rect 1346 17912 1376 17924
rect 2022 17912 2052 17924
rect 2214 17912 2244 17924
rect 2406 17912 2436 17924
rect 2598 17912 2628 17924
rect 2790 17912 2820 17924
rect 2982 17912 3012 17924
rect 3174 17912 3204 17924
rect 3850 17912 3880 17924
rect 4042 17912 4072 17924
rect 4234 17912 4264 17924
rect 4426 17912 4456 17924
rect 4618 17912 4648 17924
rect 4810 17912 4840 17924
rect 5002 17912 5032 17924
rect 5678 17912 5708 17924
rect 5870 17912 5900 17924
rect 6062 17912 6092 17924
rect 6254 17912 6284 17924
rect 6446 17912 6476 17924
rect 6638 17912 6668 17924
rect 6830 17912 6860 17924
rect 7506 17912 7536 17924
rect 7698 17912 7728 17924
rect 7890 17912 7920 17924
rect 8082 17912 8112 17924
rect 8274 17912 8304 17924
rect 8466 17912 8496 17924
rect 8658 17912 8688 17924
rect 9334 17912 9364 17924
rect 9526 17912 9556 17924
rect 9718 17912 9748 17924
rect 9910 17912 9940 17924
rect 10102 17912 10132 17924
rect 10294 17912 10324 17924
rect 10486 17912 10516 17924
rect 11162 17912 11192 17924
rect 11354 17912 11384 17924
rect 11546 17912 11576 17924
rect 11738 17912 11768 17924
rect 11930 17912 11960 17924
rect 12122 17912 12152 17924
rect 12314 17912 12344 17924
rect 12990 17912 13020 17924
rect 13182 17912 13212 17924
rect 13374 17912 13404 17924
rect 13566 17912 13596 17924
rect 13758 17912 13788 17924
rect 13950 17912 13980 17924
rect 14142 17912 14172 17924
rect 14818 17912 14848 17924
rect 15010 17912 15040 17924
rect 15202 17912 15232 17924
rect 15394 17912 15424 17924
rect 15586 17912 15616 17924
rect 15778 17912 15808 17924
rect 15970 17912 16000 17924
rect 16646 17912 16676 17924
rect 16838 17912 16868 17924
rect 17030 17912 17060 17924
rect 17222 17912 17252 17924
rect 17414 17912 17444 17924
rect 17606 17912 17636 17924
rect 17798 17912 17828 17924
rect 18474 17912 18504 17924
rect 18666 17912 18696 17924
rect 18858 17912 18888 17924
rect 19050 17912 19080 17924
rect 19242 17912 19272 17924
rect 19434 17912 19464 17924
rect 19626 17912 19656 17924
rect 20302 17912 20332 17924
rect 20494 17912 20524 17924
rect 20686 17912 20716 17924
rect 20878 17912 20908 17924
rect 21070 17912 21100 17924
rect 21262 17912 21292 17924
rect 21454 17912 21484 17924
rect 0 17853 1490 17912
rect 1828 17853 3318 17912
rect 3656 17853 5146 17912
rect 5484 17853 6974 17912
rect 7312 17853 8802 17912
rect 9140 17853 10630 17912
rect 10968 17853 12458 17912
rect 12796 17853 14286 17912
rect 14624 17853 16114 17912
rect 16452 17853 17942 17912
rect 18280 17853 19770 17912
rect 20108 17853 21598 17912
rect 0 17674 1490 17733
rect 1828 17674 3318 17733
rect 3656 17674 5146 17733
rect 5484 17674 6974 17733
rect 7312 17674 8802 17733
rect 9140 17674 10630 17733
rect 10968 17674 12458 17733
rect 12796 17674 14286 17733
rect 14624 17674 16114 17733
rect 16452 17674 17942 17733
rect 18280 17674 19770 17733
rect 20108 17674 21598 17733
rect 98 17662 128 17674
rect 290 17662 320 17674
rect 482 17662 512 17674
rect 674 17662 704 17674
rect 866 17662 896 17674
rect 1058 17662 1088 17674
rect 1250 17662 1280 17674
rect 1442 17662 1472 17674
rect 1926 17662 1956 17674
rect 2118 17662 2148 17674
rect 2310 17662 2340 17674
rect 2502 17662 2532 17674
rect 2694 17662 2724 17674
rect 2886 17662 2916 17674
rect 3078 17662 3108 17674
rect 3270 17662 3300 17674
rect 3754 17662 3784 17674
rect 3946 17662 3976 17674
rect 4138 17662 4168 17674
rect 4330 17662 4360 17674
rect 4522 17662 4552 17674
rect 4714 17662 4744 17674
rect 4906 17662 4936 17674
rect 5098 17662 5128 17674
rect 5582 17662 5612 17674
rect 5774 17662 5804 17674
rect 5966 17662 5996 17674
rect 6158 17662 6188 17674
rect 6350 17662 6380 17674
rect 6542 17662 6572 17674
rect 6734 17662 6764 17674
rect 6926 17662 6956 17674
rect 7410 17662 7440 17674
rect 7602 17662 7632 17674
rect 7794 17662 7824 17674
rect 7986 17662 8016 17674
rect 8178 17662 8208 17674
rect 8370 17662 8400 17674
rect 8562 17662 8592 17674
rect 8754 17662 8784 17674
rect 9238 17662 9268 17674
rect 9430 17662 9460 17674
rect 9622 17662 9652 17674
rect 9814 17662 9844 17674
rect 10006 17662 10036 17674
rect 10198 17662 10228 17674
rect 10390 17662 10420 17674
rect 10582 17662 10612 17674
rect 11066 17662 11096 17674
rect 11258 17662 11288 17674
rect 11450 17662 11480 17674
rect 11642 17662 11672 17674
rect 11834 17662 11864 17674
rect 12026 17662 12056 17674
rect 12218 17662 12248 17674
rect 12410 17662 12440 17674
rect 12894 17662 12924 17674
rect 13086 17662 13116 17674
rect 13278 17662 13308 17674
rect 13470 17662 13500 17674
rect 13662 17662 13692 17674
rect 13854 17662 13884 17674
rect 14046 17662 14076 17674
rect 14238 17662 14268 17674
rect 14722 17662 14752 17674
rect 14914 17662 14944 17674
rect 15106 17662 15136 17674
rect 15298 17662 15328 17674
rect 15490 17662 15520 17674
rect 15682 17662 15712 17674
rect 15874 17662 15904 17674
rect 16066 17662 16096 17674
rect 16550 17662 16580 17674
rect 16742 17662 16772 17674
rect 16934 17662 16964 17674
rect 17126 17662 17156 17674
rect 17318 17662 17348 17674
rect 17510 17662 17540 17674
rect 17702 17662 17732 17674
rect 17894 17662 17924 17674
rect 18378 17662 18408 17674
rect 18570 17662 18600 17674
rect 18762 17662 18792 17674
rect 18954 17662 18984 17674
rect 19146 17662 19176 17674
rect 19338 17662 19368 17674
rect 19530 17662 19560 17674
rect 19722 17662 19752 17674
rect 20206 17662 20236 17674
rect 20398 17662 20428 17674
rect 20590 17662 20620 17674
rect 20782 17662 20812 17674
rect 20974 17662 21004 17674
rect 21166 17662 21196 17674
rect 21358 17662 21388 17674
rect 21550 17662 21580 17674
rect 194 17198 224 17210
rect 386 17198 416 17210
rect 578 17198 608 17210
rect 770 17198 800 17210
rect 962 17198 992 17210
rect 1154 17198 1184 17210
rect 1346 17198 1376 17210
rect 2022 17198 2052 17210
rect 2214 17198 2244 17210
rect 2406 17198 2436 17210
rect 2598 17198 2628 17210
rect 2790 17198 2820 17210
rect 2982 17198 3012 17210
rect 3174 17198 3204 17210
rect 3850 17198 3880 17210
rect 4042 17198 4072 17210
rect 4234 17198 4264 17210
rect 4426 17198 4456 17210
rect 4618 17198 4648 17210
rect 4810 17198 4840 17210
rect 5002 17198 5032 17210
rect 5678 17198 5708 17210
rect 5870 17198 5900 17210
rect 6062 17198 6092 17210
rect 6254 17198 6284 17210
rect 6446 17198 6476 17210
rect 6638 17198 6668 17210
rect 6830 17198 6860 17210
rect 7506 17198 7536 17210
rect 7698 17198 7728 17210
rect 7890 17198 7920 17210
rect 8082 17198 8112 17210
rect 8274 17198 8304 17210
rect 8466 17198 8496 17210
rect 8658 17198 8688 17210
rect 9334 17198 9364 17210
rect 9526 17198 9556 17210
rect 9718 17198 9748 17210
rect 9910 17198 9940 17210
rect 10102 17198 10132 17210
rect 10294 17198 10324 17210
rect 10486 17198 10516 17210
rect 11162 17198 11192 17210
rect 11354 17198 11384 17210
rect 11546 17198 11576 17210
rect 11738 17198 11768 17210
rect 11930 17198 11960 17210
rect 12122 17198 12152 17210
rect 12314 17198 12344 17210
rect 12990 17198 13020 17210
rect 13182 17198 13212 17210
rect 13374 17198 13404 17210
rect 13566 17198 13596 17210
rect 13758 17198 13788 17210
rect 13950 17198 13980 17210
rect 14142 17198 14172 17210
rect 14818 17198 14848 17210
rect 15010 17198 15040 17210
rect 15202 17198 15232 17210
rect 15394 17198 15424 17210
rect 15586 17198 15616 17210
rect 15778 17198 15808 17210
rect 15970 17198 16000 17210
rect 16646 17198 16676 17210
rect 16838 17198 16868 17210
rect 17030 17198 17060 17210
rect 17222 17198 17252 17210
rect 17414 17198 17444 17210
rect 17606 17198 17636 17210
rect 17798 17198 17828 17210
rect 18474 17198 18504 17210
rect 18666 17198 18696 17210
rect 18858 17198 18888 17210
rect 19050 17198 19080 17210
rect 19242 17198 19272 17210
rect 19434 17198 19464 17210
rect 19626 17198 19656 17210
rect 20302 17198 20332 17210
rect 20494 17198 20524 17210
rect 20686 17198 20716 17210
rect 20878 17198 20908 17210
rect 21070 17198 21100 17210
rect 21262 17198 21292 17210
rect 21454 17198 21484 17210
rect 0 17139 1490 17198
rect 1828 17139 3318 17198
rect 3656 17139 5146 17198
rect 5484 17139 6974 17198
rect 7312 17139 8802 17198
rect 9140 17139 10630 17198
rect 10968 17139 12458 17198
rect 12796 17139 14286 17198
rect 14624 17139 16114 17198
rect 16452 17139 17942 17198
rect 18280 17139 19770 17198
rect 20108 17139 21598 17198
rect 0 16960 1490 17019
rect 1828 16960 3318 17019
rect 3656 16960 5146 17019
rect 5484 16960 6974 17019
rect 7312 16960 8802 17019
rect 9140 16960 10630 17019
rect 10968 16960 12458 17019
rect 12796 16960 14286 17019
rect 14624 16960 16114 17019
rect 16452 16960 17942 17019
rect 18280 16960 19770 17019
rect 20108 16960 21598 17019
rect 98 16948 128 16960
rect 290 16948 320 16960
rect 482 16948 512 16960
rect 674 16948 704 16960
rect 866 16948 896 16960
rect 1058 16948 1088 16960
rect 1250 16948 1280 16960
rect 1442 16948 1472 16960
rect 1926 16948 1956 16960
rect 2118 16948 2148 16960
rect 2310 16948 2340 16960
rect 2502 16948 2532 16960
rect 2694 16948 2724 16960
rect 2886 16948 2916 16960
rect 3078 16948 3108 16960
rect 3270 16948 3300 16960
rect 3754 16948 3784 16960
rect 3946 16948 3976 16960
rect 4138 16948 4168 16960
rect 4330 16948 4360 16960
rect 4522 16948 4552 16960
rect 4714 16948 4744 16960
rect 4906 16948 4936 16960
rect 5098 16948 5128 16960
rect 5582 16948 5612 16960
rect 5774 16948 5804 16960
rect 5966 16948 5996 16960
rect 6158 16948 6188 16960
rect 6350 16948 6380 16960
rect 6542 16948 6572 16960
rect 6734 16948 6764 16960
rect 6926 16948 6956 16960
rect 7410 16948 7440 16960
rect 7602 16948 7632 16960
rect 7794 16948 7824 16960
rect 7986 16948 8016 16960
rect 8178 16948 8208 16960
rect 8370 16948 8400 16960
rect 8562 16948 8592 16960
rect 8754 16948 8784 16960
rect 9238 16948 9268 16960
rect 9430 16948 9460 16960
rect 9622 16948 9652 16960
rect 9814 16948 9844 16960
rect 10006 16948 10036 16960
rect 10198 16948 10228 16960
rect 10390 16948 10420 16960
rect 10582 16948 10612 16960
rect 11066 16948 11096 16960
rect 11258 16948 11288 16960
rect 11450 16948 11480 16960
rect 11642 16948 11672 16960
rect 11834 16948 11864 16960
rect 12026 16948 12056 16960
rect 12218 16948 12248 16960
rect 12410 16948 12440 16960
rect 12894 16948 12924 16960
rect 13086 16948 13116 16960
rect 13278 16948 13308 16960
rect 13470 16948 13500 16960
rect 13662 16948 13692 16960
rect 13854 16948 13884 16960
rect 14046 16948 14076 16960
rect 14238 16948 14268 16960
rect 14722 16948 14752 16960
rect 14914 16948 14944 16960
rect 15106 16948 15136 16960
rect 15298 16948 15328 16960
rect 15490 16948 15520 16960
rect 15682 16948 15712 16960
rect 15874 16948 15904 16960
rect 16066 16948 16096 16960
rect 16550 16948 16580 16960
rect 16742 16948 16772 16960
rect 16934 16948 16964 16960
rect 17126 16948 17156 16960
rect 17318 16948 17348 16960
rect 17510 16948 17540 16960
rect 17702 16948 17732 16960
rect 17894 16948 17924 16960
rect 18378 16948 18408 16960
rect 18570 16948 18600 16960
rect 18762 16948 18792 16960
rect 18954 16948 18984 16960
rect 19146 16948 19176 16960
rect 19338 16948 19368 16960
rect 19530 16948 19560 16960
rect 19722 16948 19752 16960
rect 20206 16948 20236 16960
rect 20398 16948 20428 16960
rect 20590 16948 20620 16960
rect 20782 16948 20812 16960
rect 20974 16948 21004 16960
rect 21166 16948 21196 16960
rect 21358 16948 21388 16960
rect 21550 16948 21580 16960
rect 194 16484 224 16496
rect 386 16484 416 16496
rect 578 16484 608 16496
rect 770 16484 800 16496
rect 962 16484 992 16496
rect 1154 16484 1184 16496
rect 1346 16484 1376 16496
rect 2022 16484 2052 16496
rect 2214 16484 2244 16496
rect 2406 16484 2436 16496
rect 2598 16484 2628 16496
rect 2790 16484 2820 16496
rect 2982 16484 3012 16496
rect 3174 16484 3204 16496
rect 3850 16484 3880 16496
rect 4042 16484 4072 16496
rect 4234 16484 4264 16496
rect 4426 16484 4456 16496
rect 4618 16484 4648 16496
rect 4810 16484 4840 16496
rect 5002 16484 5032 16496
rect 5678 16484 5708 16496
rect 5870 16484 5900 16496
rect 6062 16484 6092 16496
rect 6254 16484 6284 16496
rect 6446 16484 6476 16496
rect 6638 16484 6668 16496
rect 6830 16484 6860 16496
rect 7506 16484 7536 16496
rect 7698 16484 7728 16496
rect 7890 16484 7920 16496
rect 8082 16484 8112 16496
rect 8274 16484 8304 16496
rect 8466 16484 8496 16496
rect 8658 16484 8688 16496
rect 9334 16484 9364 16496
rect 9526 16484 9556 16496
rect 9718 16484 9748 16496
rect 9910 16484 9940 16496
rect 10102 16484 10132 16496
rect 10294 16484 10324 16496
rect 10486 16484 10516 16496
rect 11162 16484 11192 16496
rect 11354 16484 11384 16496
rect 11546 16484 11576 16496
rect 11738 16484 11768 16496
rect 11930 16484 11960 16496
rect 12122 16484 12152 16496
rect 12314 16484 12344 16496
rect 12990 16484 13020 16496
rect 13182 16484 13212 16496
rect 13374 16484 13404 16496
rect 13566 16484 13596 16496
rect 13758 16484 13788 16496
rect 13950 16484 13980 16496
rect 14142 16484 14172 16496
rect 14818 16484 14848 16496
rect 15010 16484 15040 16496
rect 15202 16484 15232 16496
rect 15394 16484 15424 16496
rect 15586 16484 15616 16496
rect 15778 16484 15808 16496
rect 15970 16484 16000 16496
rect 16646 16484 16676 16496
rect 16838 16484 16868 16496
rect 17030 16484 17060 16496
rect 17222 16484 17252 16496
rect 17414 16484 17444 16496
rect 17606 16484 17636 16496
rect 17798 16484 17828 16496
rect 18474 16484 18504 16496
rect 18666 16484 18696 16496
rect 18858 16484 18888 16496
rect 19050 16484 19080 16496
rect 19242 16484 19272 16496
rect 19434 16484 19464 16496
rect 19626 16484 19656 16496
rect 20302 16484 20332 16496
rect 20494 16484 20524 16496
rect 20686 16484 20716 16496
rect 20878 16484 20908 16496
rect 21070 16484 21100 16496
rect 21262 16484 21292 16496
rect 21454 16484 21484 16496
rect 0 16425 1490 16484
rect 1828 16425 3318 16484
rect 3656 16425 5146 16484
rect 5484 16425 6974 16484
rect 7312 16425 8802 16484
rect 9140 16425 10630 16484
rect 10968 16425 12458 16484
rect 12796 16425 14286 16484
rect 14624 16425 16114 16484
rect 16452 16425 17942 16484
rect 18280 16425 19770 16484
rect 20108 16425 21598 16484
rect 0 16246 1490 16305
rect 1828 16246 3318 16305
rect 3656 16246 5146 16305
rect 5484 16246 6974 16305
rect 7312 16246 8802 16305
rect 9140 16246 10630 16305
rect 10968 16246 12458 16305
rect 12796 16246 14286 16305
rect 14624 16246 16114 16305
rect 16452 16246 17942 16305
rect 18280 16246 19770 16305
rect 20108 16246 21598 16305
rect 98 16234 128 16246
rect 290 16234 320 16246
rect 482 16234 512 16246
rect 674 16234 704 16246
rect 866 16234 896 16246
rect 1058 16234 1088 16246
rect 1250 16234 1280 16246
rect 1442 16234 1472 16246
rect 1926 16234 1956 16246
rect 2118 16234 2148 16246
rect 2310 16234 2340 16246
rect 2502 16234 2532 16246
rect 2694 16234 2724 16246
rect 2886 16234 2916 16246
rect 3078 16234 3108 16246
rect 3270 16234 3300 16246
rect 3754 16234 3784 16246
rect 3946 16234 3976 16246
rect 4138 16234 4168 16246
rect 4330 16234 4360 16246
rect 4522 16234 4552 16246
rect 4714 16234 4744 16246
rect 4906 16234 4936 16246
rect 5098 16234 5128 16246
rect 5582 16234 5612 16246
rect 5774 16234 5804 16246
rect 5966 16234 5996 16246
rect 6158 16234 6188 16246
rect 6350 16234 6380 16246
rect 6542 16234 6572 16246
rect 6734 16234 6764 16246
rect 6926 16234 6956 16246
rect 7410 16234 7440 16246
rect 7602 16234 7632 16246
rect 7794 16234 7824 16246
rect 7986 16234 8016 16246
rect 8178 16234 8208 16246
rect 8370 16234 8400 16246
rect 8562 16234 8592 16246
rect 8754 16234 8784 16246
rect 9238 16234 9268 16246
rect 9430 16234 9460 16246
rect 9622 16234 9652 16246
rect 9814 16234 9844 16246
rect 10006 16234 10036 16246
rect 10198 16234 10228 16246
rect 10390 16234 10420 16246
rect 10582 16234 10612 16246
rect 11066 16234 11096 16246
rect 11258 16234 11288 16246
rect 11450 16234 11480 16246
rect 11642 16234 11672 16246
rect 11834 16234 11864 16246
rect 12026 16234 12056 16246
rect 12218 16234 12248 16246
rect 12410 16234 12440 16246
rect 12894 16234 12924 16246
rect 13086 16234 13116 16246
rect 13278 16234 13308 16246
rect 13470 16234 13500 16246
rect 13662 16234 13692 16246
rect 13854 16234 13884 16246
rect 14046 16234 14076 16246
rect 14238 16234 14268 16246
rect 14722 16234 14752 16246
rect 14914 16234 14944 16246
rect 15106 16234 15136 16246
rect 15298 16234 15328 16246
rect 15490 16234 15520 16246
rect 15682 16234 15712 16246
rect 15874 16234 15904 16246
rect 16066 16234 16096 16246
rect 16550 16234 16580 16246
rect 16742 16234 16772 16246
rect 16934 16234 16964 16246
rect 17126 16234 17156 16246
rect 17318 16234 17348 16246
rect 17510 16234 17540 16246
rect 17702 16234 17732 16246
rect 17894 16234 17924 16246
rect 18378 16234 18408 16246
rect 18570 16234 18600 16246
rect 18762 16234 18792 16246
rect 18954 16234 18984 16246
rect 19146 16234 19176 16246
rect 19338 16234 19368 16246
rect 19530 16234 19560 16246
rect 19722 16234 19752 16246
rect 20206 16234 20236 16246
rect 20398 16234 20428 16246
rect 20590 16234 20620 16246
rect 20782 16234 20812 16246
rect 20974 16234 21004 16246
rect 21166 16234 21196 16246
rect 21358 16234 21388 16246
rect 21550 16234 21580 16246
rect 194 15770 224 15782
rect 386 15770 416 15782
rect 578 15770 608 15782
rect 770 15770 800 15782
rect 962 15770 992 15782
rect 1154 15770 1184 15782
rect 1346 15770 1376 15782
rect 2022 15770 2052 15782
rect 2214 15770 2244 15782
rect 2406 15770 2436 15782
rect 2598 15770 2628 15782
rect 2790 15770 2820 15782
rect 2982 15770 3012 15782
rect 3174 15770 3204 15782
rect 3850 15770 3880 15782
rect 4042 15770 4072 15782
rect 4234 15770 4264 15782
rect 4426 15770 4456 15782
rect 4618 15770 4648 15782
rect 4810 15770 4840 15782
rect 5002 15770 5032 15782
rect 5678 15770 5708 15782
rect 5870 15770 5900 15782
rect 6062 15770 6092 15782
rect 6254 15770 6284 15782
rect 6446 15770 6476 15782
rect 6638 15770 6668 15782
rect 6830 15770 6860 15782
rect 7506 15770 7536 15782
rect 7698 15770 7728 15782
rect 7890 15770 7920 15782
rect 8082 15770 8112 15782
rect 8274 15770 8304 15782
rect 8466 15770 8496 15782
rect 8658 15770 8688 15782
rect 9334 15770 9364 15782
rect 9526 15770 9556 15782
rect 9718 15770 9748 15782
rect 9910 15770 9940 15782
rect 10102 15770 10132 15782
rect 10294 15770 10324 15782
rect 10486 15770 10516 15782
rect 11162 15770 11192 15782
rect 11354 15770 11384 15782
rect 11546 15770 11576 15782
rect 11738 15770 11768 15782
rect 11930 15770 11960 15782
rect 12122 15770 12152 15782
rect 12314 15770 12344 15782
rect 12990 15770 13020 15782
rect 13182 15770 13212 15782
rect 13374 15770 13404 15782
rect 13566 15770 13596 15782
rect 13758 15770 13788 15782
rect 13950 15770 13980 15782
rect 14142 15770 14172 15782
rect 14818 15770 14848 15782
rect 15010 15770 15040 15782
rect 15202 15770 15232 15782
rect 15394 15770 15424 15782
rect 15586 15770 15616 15782
rect 15778 15770 15808 15782
rect 15970 15770 16000 15782
rect 16646 15770 16676 15782
rect 16838 15770 16868 15782
rect 17030 15770 17060 15782
rect 17222 15770 17252 15782
rect 17414 15770 17444 15782
rect 17606 15770 17636 15782
rect 17798 15770 17828 15782
rect 18474 15770 18504 15782
rect 18666 15770 18696 15782
rect 18858 15770 18888 15782
rect 19050 15770 19080 15782
rect 19242 15770 19272 15782
rect 19434 15770 19464 15782
rect 19626 15770 19656 15782
rect 20302 15770 20332 15782
rect 20494 15770 20524 15782
rect 20686 15770 20716 15782
rect 20878 15770 20908 15782
rect 21070 15770 21100 15782
rect 21262 15770 21292 15782
rect 21454 15770 21484 15782
rect 0 15711 1490 15770
rect 1828 15711 3318 15770
rect 3656 15711 5146 15770
rect 5484 15711 6974 15770
rect 7312 15711 8802 15770
rect 9140 15711 10630 15770
rect 10968 15711 12458 15770
rect 12796 15711 14286 15770
rect 14624 15711 16114 15770
rect 16452 15711 17942 15770
rect 18280 15711 19770 15770
rect 20108 15711 21598 15770
rect 0 15532 1490 15591
rect 1828 15532 3318 15591
rect 3656 15532 5146 15591
rect 5484 15532 6974 15591
rect 7312 15532 8802 15591
rect 9140 15532 10630 15591
rect 10968 15532 12458 15591
rect 12796 15532 14286 15591
rect 14624 15532 16114 15591
rect 16452 15532 17942 15591
rect 18280 15532 19770 15591
rect 20108 15532 21598 15591
rect 98 15520 128 15532
rect 290 15520 320 15532
rect 482 15520 512 15532
rect 674 15520 704 15532
rect 866 15520 896 15532
rect 1058 15520 1088 15532
rect 1250 15520 1280 15532
rect 1442 15520 1472 15532
rect 1926 15520 1956 15532
rect 2118 15520 2148 15532
rect 2310 15520 2340 15532
rect 2502 15520 2532 15532
rect 2694 15520 2724 15532
rect 2886 15520 2916 15532
rect 3078 15520 3108 15532
rect 3270 15520 3300 15532
rect 3754 15520 3784 15532
rect 3946 15520 3976 15532
rect 4138 15520 4168 15532
rect 4330 15520 4360 15532
rect 4522 15520 4552 15532
rect 4714 15520 4744 15532
rect 4906 15520 4936 15532
rect 5098 15520 5128 15532
rect 5582 15520 5612 15532
rect 5774 15520 5804 15532
rect 5966 15520 5996 15532
rect 6158 15520 6188 15532
rect 6350 15520 6380 15532
rect 6542 15520 6572 15532
rect 6734 15520 6764 15532
rect 6926 15520 6956 15532
rect 7410 15520 7440 15532
rect 7602 15520 7632 15532
rect 7794 15520 7824 15532
rect 7986 15520 8016 15532
rect 8178 15520 8208 15532
rect 8370 15520 8400 15532
rect 8562 15520 8592 15532
rect 8754 15520 8784 15532
rect 9238 15520 9268 15532
rect 9430 15520 9460 15532
rect 9622 15520 9652 15532
rect 9814 15520 9844 15532
rect 10006 15520 10036 15532
rect 10198 15520 10228 15532
rect 10390 15520 10420 15532
rect 10582 15520 10612 15532
rect 11066 15520 11096 15532
rect 11258 15520 11288 15532
rect 11450 15520 11480 15532
rect 11642 15520 11672 15532
rect 11834 15520 11864 15532
rect 12026 15520 12056 15532
rect 12218 15520 12248 15532
rect 12410 15520 12440 15532
rect 12894 15520 12924 15532
rect 13086 15520 13116 15532
rect 13278 15520 13308 15532
rect 13470 15520 13500 15532
rect 13662 15520 13692 15532
rect 13854 15520 13884 15532
rect 14046 15520 14076 15532
rect 14238 15520 14268 15532
rect 14722 15520 14752 15532
rect 14914 15520 14944 15532
rect 15106 15520 15136 15532
rect 15298 15520 15328 15532
rect 15490 15520 15520 15532
rect 15682 15520 15712 15532
rect 15874 15520 15904 15532
rect 16066 15520 16096 15532
rect 16550 15520 16580 15532
rect 16742 15520 16772 15532
rect 16934 15520 16964 15532
rect 17126 15520 17156 15532
rect 17318 15520 17348 15532
rect 17510 15520 17540 15532
rect 17702 15520 17732 15532
rect 17894 15520 17924 15532
rect 18378 15520 18408 15532
rect 18570 15520 18600 15532
rect 18762 15520 18792 15532
rect 18954 15520 18984 15532
rect 19146 15520 19176 15532
rect 19338 15520 19368 15532
rect 19530 15520 19560 15532
rect 19722 15520 19752 15532
rect 20206 15520 20236 15532
rect 20398 15520 20428 15532
rect 20590 15520 20620 15532
rect 20782 15520 20812 15532
rect 20974 15520 21004 15532
rect 21166 15520 21196 15532
rect 21358 15520 21388 15532
rect 21550 15520 21580 15532
rect 194 15056 224 15068
rect 386 15056 416 15068
rect 578 15056 608 15068
rect 770 15056 800 15068
rect 962 15056 992 15068
rect 1154 15056 1184 15068
rect 1346 15056 1376 15068
rect 2022 15056 2052 15068
rect 2214 15056 2244 15068
rect 2406 15056 2436 15068
rect 2598 15056 2628 15068
rect 2790 15056 2820 15068
rect 2982 15056 3012 15068
rect 3174 15056 3204 15068
rect 3850 15056 3880 15068
rect 4042 15056 4072 15068
rect 4234 15056 4264 15068
rect 4426 15056 4456 15068
rect 4618 15056 4648 15068
rect 4810 15056 4840 15068
rect 5002 15056 5032 15068
rect 5678 15056 5708 15068
rect 5870 15056 5900 15068
rect 6062 15056 6092 15068
rect 6254 15056 6284 15068
rect 6446 15056 6476 15068
rect 6638 15056 6668 15068
rect 6830 15056 6860 15068
rect 7506 15056 7536 15068
rect 7698 15056 7728 15068
rect 7890 15056 7920 15068
rect 8082 15056 8112 15068
rect 8274 15056 8304 15068
rect 8466 15056 8496 15068
rect 8658 15056 8688 15068
rect 9334 15056 9364 15068
rect 9526 15056 9556 15068
rect 9718 15056 9748 15068
rect 9910 15056 9940 15068
rect 10102 15056 10132 15068
rect 10294 15056 10324 15068
rect 10486 15056 10516 15068
rect 11162 15056 11192 15068
rect 11354 15056 11384 15068
rect 11546 15056 11576 15068
rect 11738 15056 11768 15068
rect 11930 15056 11960 15068
rect 12122 15056 12152 15068
rect 12314 15056 12344 15068
rect 12990 15056 13020 15068
rect 13182 15056 13212 15068
rect 13374 15056 13404 15068
rect 13566 15056 13596 15068
rect 13758 15056 13788 15068
rect 13950 15056 13980 15068
rect 14142 15056 14172 15068
rect 14818 15056 14848 15068
rect 15010 15056 15040 15068
rect 15202 15056 15232 15068
rect 15394 15056 15424 15068
rect 15586 15056 15616 15068
rect 15778 15056 15808 15068
rect 15970 15056 16000 15068
rect 16646 15056 16676 15068
rect 16838 15056 16868 15068
rect 17030 15056 17060 15068
rect 17222 15056 17252 15068
rect 17414 15056 17444 15068
rect 17606 15056 17636 15068
rect 17798 15056 17828 15068
rect 18474 15056 18504 15068
rect 18666 15056 18696 15068
rect 18858 15056 18888 15068
rect 19050 15056 19080 15068
rect 19242 15056 19272 15068
rect 19434 15056 19464 15068
rect 19626 15056 19656 15068
rect 20302 15056 20332 15068
rect 20494 15056 20524 15068
rect 20686 15056 20716 15068
rect 20878 15056 20908 15068
rect 21070 15056 21100 15068
rect 21262 15056 21292 15068
rect 21454 15056 21484 15068
rect 0 14997 1490 15056
rect 1828 14997 3318 15056
rect 3656 14997 5146 15056
rect 5484 14997 6974 15056
rect 7312 14997 8802 15056
rect 9140 14997 10630 15056
rect 10968 14997 12458 15056
rect 12796 14997 14286 15056
rect 14624 14997 16114 15056
rect 16452 14997 17942 15056
rect 18280 14997 19770 15056
rect 20108 14997 21598 15056
rect 0 14818 1490 14877
rect 1828 14818 3318 14877
rect 3656 14818 5146 14877
rect 5484 14818 6974 14877
rect 7312 14818 8802 14877
rect 9140 14818 10630 14877
rect 10968 14818 12458 14877
rect 12796 14818 14286 14877
rect 14624 14818 16114 14877
rect 16452 14818 17942 14877
rect 18280 14818 19770 14877
rect 20108 14818 21598 14877
rect 98 14806 128 14818
rect 290 14806 320 14818
rect 482 14806 512 14818
rect 674 14806 704 14818
rect 866 14806 896 14818
rect 1058 14806 1088 14818
rect 1250 14806 1280 14818
rect 1442 14806 1472 14818
rect 1926 14806 1956 14818
rect 2118 14806 2148 14818
rect 2310 14806 2340 14818
rect 2502 14806 2532 14818
rect 2694 14806 2724 14818
rect 2886 14806 2916 14818
rect 3078 14806 3108 14818
rect 3270 14806 3300 14818
rect 3754 14806 3784 14818
rect 3946 14806 3976 14818
rect 4138 14806 4168 14818
rect 4330 14806 4360 14818
rect 4522 14806 4552 14818
rect 4714 14806 4744 14818
rect 4906 14806 4936 14818
rect 5098 14806 5128 14818
rect 5582 14806 5612 14818
rect 5774 14806 5804 14818
rect 5966 14806 5996 14818
rect 6158 14806 6188 14818
rect 6350 14806 6380 14818
rect 6542 14806 6572 14818
rect 6734 14806 6764 14818
rect 6926 14806 6956 14818
rect 7410 14806 7440 14818
rect 7602 14806 7632 14818
rect 7794 14806 7824 14818
rect 7986 14806 8016 14818
rect 8178 14806 8208 14818
rect 8370 14806 8400 14818
rect 8562 14806 8592 14818
rect 8754 14806 8784 14818
rect 9238 14806 9268 14818
rect 9430 14806 9460 14818
rect 9622 14806 9652 14818
rect 9814 14806 9844 14818
rect 10006 14806 10036 14818
rect 10198 14806 10228 14818
rect 10390 14806 10420 14818
rect 10582 14806 10612 14818
rect 11066 14806 11096 14818
rect 11258 14806 11288 14818
rect 11450 14806 11480 14818
rect 11642 14806 11672 14818
rect 11834 14806 11864 14818
rect 12026 14806 12056 14818
rect 12218 14806 12248 14818
rect 12410 14806 12440 14818
rect 12894 14806 12924 14818
rect 13086 14806 13116 14818
rect 13278 14806 13308 14818
rect 13470 14806 13500 14818
rect 13662 14806 13692 14818
rect 13854 14806 13884 14818
rect 14046 14806 14076 14818
rect 14238 14806 14268 14818
rect 14722 14806 14752 14818
rect 14914 14806 14944 14818
rect 15106 14806 15136 14818
rect 15298 14806 15328 14818
rect 15490 14806 15520 14818
rect 15682 14806 15712 14818
rect 15874 14806 15904 14818
rect 16066 14806 16096 14818
rect 16550 14806 16580 14818
rect 16742 14806 16772 14818
rect 16934 14806 16964 14818
rect 17126 14806 17156 14818
rect 17318 14806 17348 14818
rect 17510 14806 17540 14818
rect 17702 14806 17732 14818
rect 17894 14806 17924 14818
rect 18378 14806 18408 14818
rect 18570 14806 18600 14818
rect 18762 14806 18792 14818
rect 18954 14806 18984 14818
rect 19146 14806 19176 14818
rect 19338 14806 19368 14818
rect 19530 14806 19560 14818
rect 19722 14806 19752 14818
rect 20206 14806 20236 14818
rect 20398 14806 20428 14818
rect 20590 14806 20620 14818
rect 20782 14806 20812 14818
rect 20974 14806 21004 14818
rect 21166 14806 21196 14818
rect 21358 14806 21388 14818
rect 21550 14806 21580 14818
rect 194 14342 224 14354
rect 386 14342 416 14354
rect 578 14342 608 14354
rect 770 14342 800 14354
rect 962 14342 992 14354
rect 1154 14342 1184 14354
rect 1346 14342 1376 14354
rect 2022 14342 2052 14354
rect 2214 14342 2244 14354
rect 2406 14342 2436 14354
rect 2598 14342 2628 14354
rect 2790 14342 2820 14354
rect 2982 14342 3012 14354
rect 3174 14342 3204 14354
rect 3850 14342 3880 14354
rect 4042 14342 4072 14354
rect 4234 14342 4264 14354
rect 4426 14342 4456 14354
rect 4618 14342 4648 14354
rect 4810 14342 4840 14354
rect 5002 14342 5032 14354
rect 5678 14342 5708 14354
rect 5870 14342 5900 14354
rect 6062 14342 6092 14354
rect 6254 14342 6284 14354
rect 6446 14342 6476 14354
rect 6638 14342 6668 14354
rect 6830 14342 6860 14354
rect 7506 14342 7536 14354
rect 7698 14342 7728 14354
rect 7890 14342 7920 14354
rect 8082 14342 8112 14354
rect 8274 14342 8304 14354
rect 8466 14342 8496 14354
rect 8658 14342 8688 14354
rect 9334 14342 9364 14354
rect 9526 14342 9556 14354
rect 9718 14342 9748 14354
rect 9910 14342 9940 14354
rect 10102 14342 10132 14354
rect 10294 14342 10324 14354
rect 10486 14342 10516 14354
rect 11162 14342 11192 14354
rect 11354 14342 11384 14354
rect 11546 14342 11576 14354
rect 11738 14342 11768 14354
rect 11930 14342 11960 14354
rect 12122 14342 12152 14354
rect 12314 14342 12344 14354
rect 12990 14342 13020 14354
rect 13182 14342 13212 14354
rect 13374 14342 13404 14354
rect 13566 14342 13596 14354
rect 13758 14342 13788 14354
rect 13950 14342 13980 14354
rect 14142 14342 14172 14354
rect 14818 14342 14848 14354
rect 15010 14342 15040 14354
rect 15202 14342 15232 14354
rect 15394 14342 15424 14354
rect 15586 14342 15616 14354
rect 15778 14342 15808 14354
rect 15970 14342 16000 14354
rect 16646 14342 16676 14354
rect 16838 14342 16868 14354
rect 17030 14342 17060 14354
rect 17222 14342 17252 14354
rect 17414 14342 17444 14354
rect 17606 14342 17636 14354
rect 17798 14342 17828 14354
rect 18474 14342 18504 14354
rect 18666 14342 18696 14354
rect 18858 14342 18888 14354
rect 19050 14342 19080 14354
rect 19242 14342 19272 14354
rect 19434 14342 19464 14354
rect 19626 14342 19656 14354
rect 20302 14342 20332 14354
rect 20494 14342 20524 14354
rect 20686 14342 20716 14354
rect 20878 14342 20908 14354
rect 21070 14342 21100 14354
rect 21262 14342 21292 14354
rect 21454 14342 21484 14354
rect 0 14283 1490 14342
rect 1828 14283 3318 14342
rect 3656 14283 5146 14342
rect 5484 14283 6974 14342
rect 7312 14283 8802 14342
rect 9140 14283 10630 14342
rect 10968 14283 12458 14342
rect 12796 14283 14286 14342
rect 14624 14283 16114 14342
rect 16452 14283 17942 14342
rect 18280 14283 19770 14342
rect 20108 14283 21598 14342
rect 0 14104 1490 14163
rect 1828 14104 3318 14163
rect 3656 14104 5146 14163
rect 5484 14104 6974 14163
rect 7312 14104 8802 14163
rect 9140 14104 10630 14163
rect 10968 14104 12458 14163
rect 12796 14104 14286 14163
rect 14624 14104 16114 14163
rect 16452 14104 17942 14163
rect 18280 14104 19770 14163
rect 20108 14104 21598 14163
rect 98 14092 128 14104
rect 290 14092 320 14104
rect 482 14092 512 14104
rect 674 14092 704 14104
rect 866 14092 896 14104
rect 1058 14092 1088 14104
rect 1250 14092 1280 14104
rect 1442 14092 1472 14104
rect 1926 14092 1956 14104
rect 2118 14092 2148 14104
rect 2310 14092 2340 14104
rect 2502 14092 2532 14104
rect 2694 14092 2724 14104
rect 2886 14092 2916 14104
rect 3078 14092 3108 14104
rect 3270 14092 3300 14104
rect 3754 14092 3784 14104
rect 3946 14092 3976 14104
rect 4138 14092 4168 14104
rect 4330 14092 4360 14104
rect 4522 14092 4552 14104
rect 4714 14092 4744 14104
rect 4906 14092 4936 14104
rect 5098 14092 5128 14104
rect 5582 14092 5612 14104
rect 5774 14092 5804 14104
rect 5966 14092 5996 14104
rect 6158 14092 6188 14104
rect 6350 14092 6380 14104
rect 6542 14092 6572 14104
rect 6734 14092 6764 14104
rect 6926 14092 6956 14104
rect 7410 14092 7440 14104
rect 7602 14092 7632 14104
rect 7794 14092 7824 14104
rect 7986 14092 8016 14104
rect 8178 14092 8208 14104
rect 8370 14092 8400 14104
rect 8562 14092 8592 14104
rect 8754 14092 8784 14104
rect 9238 14092 9268 14104
rect 9430 14092 9460 14104
rect 9622 14092 9652 14104
rect 9814 14092 9844 14104
rect 10006 14092 10036 14104
rect 10198 14092 10228 14104
rect 10390 14092 10420 14104
rect 10582 14092 10612 14104
rect 11066 14092 11096 14104
rect 11258 14092 11288 14104
rect 11450 14092 11480 14104
rect 11642 14092 11672 14104
rect 11834 14092 11864 14104
rect 12026 14092 12056 14104
rect 12218 14092 12248 14104
rect 12410 14092 12440 14104
rect 12894 14092 12924 14104
rect 13086 14092 13116 14104
rect 13278 14092 13308 14104
rect 13470 14092 13500 14104
rect 13662 14092 13692 14104
rect 13854 14092 13884 14104
rect 14046 14092 14076 14104
rect 14238 14092 14268 14104
rect 14722 14092 14752 14104
rect 14914 14092 14944 14104
rect 15106 14092 15136 14104
rect 15298 14092 15328 14104
rect 15490 14092 15520 14104
rect 15682 14092 15712 14104
rect 15874 14092 15904 14104
rect 16066 14092 16096 14104
rect 16550 14092 16580 14104
rect 16742 14092 16772 14104
rect 16934 14092 16964 14104
rect 17126 14092 17156 14104
rect 17318 14092 17348 14104
rect 17510 14092 17540 14104
rect 17702 14092 17732 14104
rect 17894 14092 17924 14104
rect 18378 14092 18408 14104
rect 18570 14092 18600 14104
rect 18762 14092 18792 14104
rect 18954 14092 18984 14104
rect 19146 14092 19176 14104
rect 19338 14092 19368 14104
rect 19530 14092 19560 14104
rect 19722 14092 19752 14104
rect 20206 14092 20236 14104
rect 20398 14092 20428 14104
rect 20590 14092 20620 14104
rect 20782 14092 20812 14104
rect 20974 14092 21004 14104
rect 21166 14092 21196 14104
rect 21358 14092 21388 14104
rect 21550 14092 21580 14104
rect 194 13628 224 13640
rect 386 13628 416 13640
rect 578 13628 608 13640
rect 770 13628 800 13640
rect 962 13628 992 13640
rect 1154 13628 1184 13640
rect 1346 13628 1376 13640
rect 2022 13628 2052 13640
rect 2214 13628 2244 13640
rect 2406 13628 2436 13640
rect 2598 13628 2628 13640
rect 2790 13628 2820 13640
rect 2982 13628 3012 13640
rect 3174 13628 3204 13640
rect 3850 13628 3880 13640
rect 4042 13628 4072 13640
rect 4234 13628 4264 13640
rect 4426 13628 4456 13640
rect 4618 13628 4648 13640
rect 4810 13628 4840 13640
rect 5002 13628 5032 13640
rect 5678 13628 5708 13640
rect 5870 13628 5900 13640
rect 6062 13628 6092 13640
rect 6254 13628 6284 13640
rect 6446 13628 6476 13640
rect 6638 13628 6668 13640
rect 6830 13628 6860 13640
rect 7506 13628 7536 13640
rect 7698 13628 7728 13640
rect 7890 13628 7920 13640
rect 8082 13628 8112 13640
rect 8274 13628 8304 13640
rect 8466 13628 8496 13640
rect 8658 13628 8688 13640
rect 9334 13628 9364 13640
rect 9526 13628 9556 13640
rect 9718 13628 9748 13640
rect 9910 13628 9940 13640
rect 10102 13628 10132 13640
rect 10294 13628 10324 13640
rect 10486 13628 10516 13640
rect 11162 13628 11192 13640
rect 11354 13628 11384 13640
rect 11546 13628 11576 13640
rect 11738 13628 11768 13640
rect 11930 13628 11960 13640
rect 12122 13628 12152 13640
rect 12314 13628 12344 13640
rect 12990 13628 13020 13640
rect 13182 13628 13212 13640
rect 13374 13628 13404 13640
rect 13566 13628 13596 13640
rect 13758 13628 13788 13640
rect 13950 13628 13980 13640
rect 14142 13628 14172 13640
rect 14818 13628 14848 13640
rect 15010 13628 15040 13640
rect 15202 13628 15232 13640
rect 15394 13628 15424 13640
rect 15586 13628 15616 13640
rect 15778 13628 15808 13640
rect 15970 13628 16000 13640
rect 16646 13628 16676 13640
rect 16838 13628 16868 13640
rect 17030 13628 17060 13640
rect 17222 13628 17252 13640
rect 17414 13628 17444 13640
rect 17606 13628 17636 13640
rect 17798 13628 17828 13640
rect 18474 13628 18504 13640
rect 18666 13628 18696 13640
rect 18858 13628 18888 13640
rect 19050 13628 19080 13640
rect 19242 13628 19272 13640
rect 19434 13628 19464 13640
rect 19626 13628 19656 13640
rect 20302 13628 20332 13640
rect 20494 13628 20524 13640
rect 20686 13628 20716 13640
rect 20878 13628 20908 13640
rect 21070 13628 21100 13640
rect 21262 13628 21292 13640
rect 21454 13628 21484 13640
rect 0 13569 1490 13628
rect 1828 13569 3318 13628
rect 3656 13569 5146 13628
rect 5484 13569 6974 13628
rect 7312 13569 8802 13628
rect 9140 13569 10630 13628
rect 10968 13569 12458 13628
rect 12796 13569 14286 13628
rect 14624 13569 16114 13628
rect 16452 13569 17942 13628
rect 18280 13569 19770 13628
rect 20108 13569 21598 13628
rect 0 13390 1490 13449
rect 1828 13390 3318 13449
rect 3656 13390 5146 13449
rect 5484 13390 6974 13449
rect 7312 13390 8802 13449
rect 9140 13390 10630 13449
rect 10968 13390 12458 13449
rect 12796 13390 14286 13449
rect 14624 13390 16114 13449
rect 16452 13390 17942 13449
rect 18280 13390 19770 13449
rect 20108 13390 21598 13449
rect 98 13378 128 13390
rect 290 13378 320 13390
rect 482 13378 512 13390
rect 674 13378 704 13390
rect 866 13378 896 13390
rect 1058 13378 1088 13390
rect 1250 13378 1280 13390
rect 1442 13378 1472 13390
rect 1926 13378 1956 13390
rect 2118 13378 2148 13390
rect 2310 13378 2340 13390
rect 2502 13378 2532 13390
rect 2694 13378 2724 13390
rect 2886 13378 2916 13390
rect 3078 13378 3108 13390
rect 3270 13378 3300 13390
rect 3754 13378 3784 13390
rect 3946 13378 3976 13390
rect 4138 13378 4168 13390
rect 4330 13378 4360 13390
rect 4522 13378 4552 13390
rect 4714 13378 4744 13390
rect 4906 13378 4936 13390
rect 5098 13378 5128 13390
rect 5582 13378 5612 13390
rect 5774 13378 5804 13390
rect 5966 13378 5996 13390
rect 6158 13378 6188 13390
rect 6350 13378 6380 13390
rect 6542 13378 6572 13390
rect 6734 13378 6764 13390
rect 6926 13378 6956 13390
rect 7410 13378 7440 13390
rect 7602 13378 7632 13390
rect 7794 13378 7824 13390
rect 7986 13378 8016 13390
rect 8178 13378 8208 13390
rect 8370 13378 8400 13390
rect 8562 13378 8592 13390
rect 8754 13378 8784 13390
rect 9238 13378 9268 13390
rect 9430 13378 9460 13390
rect 9622 13378 9652 13390
rect 9814 13378 9844 13390
rect 10006 13378 10036 13390
rect 10198 13378 10228 13390
rect 10390 13378 10420 13390
rect 10582 13378 10612 13390
rect 11066 13378 11096 13390
rect 11258 13378 11288 13390
rect 11450 13378 11480 13390
rect 11642 13378 11672 13390
rect 11834 13378 11864 13390
rect 12026 13378 12056 13390
rect 12218 13378 12248 13390
rect 12410 13378 12440 13390
rect 12894 13378 12924 13390
rect 13086 13378 13116 13390
rect 13278 13378 13308 13390
rect 13470 13378 13500 13390
rect 13662 13378 13692 13390
rect 13854 13378 13884 13390
rect 14046 13378 14076 13390
rect 14238 13378 14268 13390
rect 14722 13378 14752 13390
rect 14914 13378 14944 13390
rect 15106 13378 15136 13390
rect 15298 13378 15328 13390
rect 15490 13378 15520 13390
rect 15682 13378 15712 13390
rect 15874 13378 15904 13390
rect 16066 13378 16096 13390
rect 16550 13378 16580 13390
rect 16742 13378 16772 13390
rect 16934 13378 16964 13390
rect 17126 13378 17156 13390
rect 17318 13378 17348 13390
rect 17510 13378 17540 13390
rect 17702 13378 17732 13390
rect 17894 13378 17924 13390
rect 18378 13378 18408 13390
rect 18570 13378 18600 13390
rect 18762 13378 18792 13390
rect 18954 13378 18984 13390
rect 19146 13378 19176 13390
rect 19338 13378 19368 13390
rect 19530 13378 19560 13390
rect 19722 13378 19752 13390
rect 20206 13378 20236 13390
rect 20398 13378 20428 13390
rect 20590 13378 20620 13390
rect 20782 13378 20812 13390
rect 20974 13378 21004 13390
rect 21166 13378 21196 13390
rect 21358 13378 21388 13390
rect 21550 13378 21580 13390
rect 194 12914 224 12926
rect 386 12914 416 12926
rect 578 12914 608 12926
rect 770 12914 800 12926
rect 962 12914 992 12926
rect 1154 12914 1184 12926
rect 1346 12914 1376 12926
rect 2022 12914 2052 12926
rect 2214 12914 2244 12926
rect 2406 12914 2436 12926
rect 2598 12914 2628 12926
rect 2790 12914 2820 12926
rect 2982 12914 3012 12926
rect 3174 12914 3204 12926
rect 3850 12914 3880 12926
rect 4042 12914 4072 12926
rect 4234 12914 4264 12926
rect 4426 12914 4456 12926
rect 4618 12914 4648 12926
rect 4810 12914 4840 12926
rect 5002 12914 5032 12926
rect 5678 12914 5708 12926
rect 5870 12914 5900 12926
rect 6062 12914 6092 12926
rect 6254 12914 6284 12926
rect 6446 12914 6476 12926
rect 6638 12914 6668 12926
rect 6830 12914 6860 12926
rect 7506 12914 7536 12926
rect 7698 12914 7728 12926
rect 7890 12914 7920 12926
rect 8082 12914 8112 12926
rect 8274 12914 8304 12926
rect 8466 12914 8496 12926
rect 8658 12914 8688 12926
rect 9334 12914 9364 12926
rect 9526 12914 9556 12926
rect 9718 12914 9748 12926
rect 9910 12914 9940 12926
rect 10102 12914 10132 12926
rect 10294 12914 10324 12926
rect 10486 12914 10516 12926
rect 11162 12914 11192 12926
rect 11354 12914 11384 12926
rect 11546 12914 11576 12926
rect 11738 12914 11768 12926
rect 11930 12914 11960 12926
rect 12122 12914 12152 12926
rect 12314 12914 12344 12926
rect 12990 12914 13020 12926
rect 13182 12914 13212 12926
rect 13374 12914 13404 12926
rect 13566 12914 13596 12926
rect 13758 12914 13788 12926
rect 13950 12914 13980 12926
rect 14142 12914 14172 12926
rect 14818 12914 14848 12926
rect 15010 12914 15040 12926
rect 15202 12914 15232 12926
rect 15394 12914 15424 12926
rect 15586 12914 15616 12926
rect 15778 12914 15808 12926
rect 15970 12914 16000 12926
rect 16646 12914 16676 12926
rect 16838 12914 16868 12926
rect 17030 12914 17060 12926
rect 17222 12914 17252 12926
rect 17414 12914 17444 12926
rect 17606 12914 17636 12926
rect 17798 12914 17828 12926
rect 18474 12914 18504 12926
rect 18666 12914 18696 12926
rect 18858 12914 18888 12926
rect 19050 12914 19080 12926
rect 19242 12914 19272 12926
rect 19434 12914 19464 12926
rect 19626 12914 19656 12926
rect 20302 12914 20332 12926
rect 20494 12914 20524 12926
rect 20686 12914 20716 12926
rect 20878 12914 20908 12926
rect 21070 12914 21100 12926
rect 21262 12914 21292 12926
rect 21454 12914 21484 12926
rect 0 12855 1490 12914
rect 1828 12855 3318 12914
rect 3656 12855 5146 12914
rect 5484 12855 6974 12914
rect 7312 12855 8802 12914
rect 9140 12855 10630 12914
rect 10968 12855 12458 12914
rect 12796 12855 14286 12914
rect 14624 12855 16114 12914
rect 16452 12855 17942 12914
rect 18280 12855 19770 12914
rect 20108 12855 21598 12914
rect 0 12676 1490 12735
rect 1828 12676 3318 12735
rect 3656 12676 5146 12735
rect 5484 12676 6974 12735
rect 7312 12676 8802 12735
rect 9140 12676 10630 12735
rect 10968 12676 12458 12735
rect 12796 12676 14286 12735
rect 14624 12676 16114 12735
rect 16452 12676 17942 12735
rect 18280 12676 19770 12735
rect 20108 12676 21598 12735
rect 98 12664 128 12676
rect 290 12664 320 12676
rect 482 12664 512 12676
rect 674 12664 704 12676
rect 866 12664 896 12676
rect 1058 12664 1088 12676
rect 1250 12664 1280 12676
rect 1442 12664 1472 12676
rect 1926 12664 1956 12676
rect 2118 12664 2148 12676
rect 2310 12664 2340 12676
rect 2502 12664 2532 12676
rect 2694 12664 2724 12676
rect 2886 12664 2916 12676
rect 3078 12664 3108 12676
rect 3270 12664 3300 12676
rect 3754 12664 3784 12676
rect 3946 12664 3976 12676
rect 4138 12664 4168 12676
rect 4330 12664 4360 12676
rect 4522 12664 4552 12676
rect 4714 12664 4744 12676
rect 4906 12664 4936 12676
rect 5098 12664 5128 12676
rect 5582 12664 5612 12676
rect 5774 12664 5804 12676
rect 5966 12664 5996 12676
rect 6158 12664 6188 12676
rect 6350 12664 6380 12676
rect 6542 12664 6572 12676
rect 6734 12664 6764 12676
rect 6926 12664 6956 12676
rect 7410 12664 7440 12676
rect 7602 12664 7632 12676
rect 7794 12664 7824 12676
rect 7986 12664 8016 12676
rect 8178 12664 8208 12676
rect 8370 12664 8400 12676
rect 8562 12664 8592 12676
rect 8754 12664 8784 12676
rect 9238 12664 9268 12676
rect 9430 12664 9460 12676
rect 9622 12664 9652 12676
rect 9814 12664 9844 12676
rect 10006 12664 10036 12676
rect 10198 12664 10228 12676
rect 10390 12664 10420 12676
rect 10582 12664 10612 12676
rect 11066 12664 11096 12676
rect 11258 12664 11288 12676
rect 11450 12664 11480 12676
rect 11642 12664 11672 12676
rect 11834 12664 11864 12676
rect 12026 12664 12056 12676
rect 12218 12664 12248 12676
rect 12410 12664 12440 12676
rect 12894 12664 12924 12676
rect 13086 12664 13116 12676
rect 13278 12664 13308 12676
rect 13470 12664 13500 12676
rect 13662 12664 13692 12676
rect 13854 12664 13884 12676
rect 14046 12664 14076 12676
rect 14238 12664 14268 12676
rect 14722 12664 14752 12676
rect 14914 12664 14944 12676
rect 15106 12664 15136 12676
rect 15298 12664 15328 12676
rect 15490 12664 15520 12676
rect 15682 12664 15712 12676
rect 15874 12664 15904 12676
rect 16066 12664 16096 12676
rect 16550 12664 16580 12676
rect 16742 12664 16772 12676
rect 16934 12664 16964 12676
rect 17126 12664 17156 12676
rect 17318 12664 17348 12676
rect 17510 12664 17540 12676
rect 17702 12664 17732 12676
rect 17894 12664 17924 12676
rect 18378 12664 18408 12676
rect 18570 12664 18600 12676
rect 18762 12664 18792 12676
rect 18954 12664 18984 12676
rect 19146 12664 19176 12676
rect 19338 12664 19368 12676
rect 19530 12664 19560 12676
rect 19722 12664 19752 12676
rect 20206 12664 20236 12676
rect 20398 12664 20428 12676
rect 20590 12664 20620 12676
rect 20782 12664 20812 12676
rect 20974 12664 21004 12676
rect 21166 12664 21196 12676
rect 21358 12664 21388 12676
rect 21550 12664 21580 12676
rect 194 12200 224 12212
rect 386 12200 416 12212
rect 578 12200 608 12212
rect 770 12200 800 12212
rect 962 12200 992 12212
rect 1154 12200 1184 12212
rect 1346 12200 1376 12212
rect 2022 12200 2052 12212
rect 2214 12200 2244 12212
rect 2406 12200 2436 12212
rect 2598 12200 2628 12212
rect 2790 12200 2820 12212
rect 2982 12200 3012 12212
rect 3174 12200 3204 12212
rect 3850 12200 3880 12212
rect 4042 12200 4072 12212
rect 4234 12200 4264 12212
rect 4426 12200 4456 12212
rect 4618 12200 4648 12212
rect 4810 12200 4840 12212
rect 5002 12200 5032 12212
rect 5678 12200 5708 12212
rect 5870 12200 5900 12212
rect 6062 12200 6092 12212
rect 6254 12200 6284 12212
rect 6446 12200 6476 12212
rect 6638 12200 6668 12212
rect 6830 12200 6860 12212
rect 7506 12200 7536 12212
rect 7698 12200 7728 12212
rect 7890 12200 7920 12212
rect 8082 12200 8112 12212
rect 8274 12200 8304 12212
rect 8466 12200 8496 12212
rect 8658 12200 8688 12212
rect 9334 12200 9364 12212
rect 9526 12200 9556 12212
rect 9718 12200 9748 12212
rect 9910 12200 9940 12212
rect 10102 12200 10132 12212
rect 10294 12200 10324 12212
rect 10486 12200 10516 12212
rect 11162 12200 11192 12212
rect 11354 12200 11384 12212
rect 11546 12200 11576 12212
rect 11738 12200 11768 12212
rect 11930 12200 11960 12212
rect 12122 12200 12152 12212
rect 12314 12200 12344 12212
rect 12990 12200 13020 12212
rect 13182 12200 13212 12212
rect 13374 12200 13404 12212
rect 13566 12200 13596 12212
rect 13758 12200 13788 12212
rect 13950 12200 13980 12212
rect 14142 12200 14172 12212
rect 14818 12200 14848 12212
rect 15010 12200 15040 12212
rect 15202 12200 15232 12212
rect 15394 12200 15424 12212
rect 15586 12200 15616 12212
rect 15778 12200 15808 12212
rect 15970 12200 16000 12212
rect 16646 12200 16676 12212
rect 16838 12200 16868 12212
rect 17030 12200 17060 12212
rect 17222 12200 17252 12212
rect 17414 12200 17444 12212
rect 17606 12200 17636 12212
rect 17798 12200 17828 12212
rect 18474 12200 18504 12212
rect 18666 12200 18696 12212
rect 18858 12200 18888 12212
rect 19050 12200 19080 12212
rect 19242 12200 19272 12212
rect 19434 12200 19464 12212
rect 19626 12200 19656 12212
rect 20302 12200 20332 12212
rect 20494 12200 20524 12212
rect 20686 12200 20716 12212
rect 20878 12200 20908 12212
rect 21070 12200 21100 12212
rect 21262 12200 21292 12212
rect 21454 12200 21484 12212
rect 0 12141 1490 12200
rect 1828 12141 3318 12200
rect 3656 12141 5146 12200
rect 5484 12141 6974 12200
rect 7312 12141 8802 12200
rect 9140 12141 10630 12200
rect 10968 12141 12458 12200
rect 12796 12141 14286 12200
rect 14624 12141 16114 12200
rect 16452 12141 17942 12200
rect 18280 12141 19770 12200
rect 20108 12141 21598 12200
rect 0 11962 1490 12021
rect 1828 11962 3318 12021
rect 3656 11962 5146 12021
rect 5484 11962 6974 12021
rect 7312 11962 8802 12021
rect 9140 11962 10630 12021
rect 10968 11962 12458 12021
rect 12796 11962 14286 12021
rect 14624 11962 16114 12021
rect 16452 11962 17942 12021
rect 18280 11962 19770 12021
rect 20108 11962 21598 12021
rect 98 11950 128 11962
rect 290 11950 320 11962
rect 482 11950 512 11962
rect 674 11950 704 11962
rect 866 11950 896 11962
rect 1058 11950 1088 11962
rect 1250 11950 1280 11962
rect 1442 11950 1472 11962
rect 1926 11950 1956 11962
rect 2118 11950 2148 11962
rect 2310 11950 2340 11962
rect 2502 11950 2532 11962
rect 2694 11950 2724 11962
rect 2886 11950 2916 11962
rect 3078 11950 3108 11962
rect 3270 11950 3300 11962
rect 3754 11950 3784 11962
rect 3946 11950 3976 11962
rect 4138 11950 4168 11962
rect 4330 11950 4360 11962
rect 4522 11950 4552 11962
rect 4714 11950 4744 11962
rect 4906 11950 4936 11962
rect 5098 11950 5128 11962
rect 5582 11950 5612 11962
rect 5774 11950 5804 11962
rect 5966 11950 5996 11962
rect 6158 11950 6188 11962
rect 6350 11950 6380 11962
rect 6542 11950 6572 11962
rect 6734 11950 6764 11962
rect 6926 11950 6956 11962
rect 7410 11950 7440 11962
rect 7602 11950 7632 11962
rect 7794 11950 7824 11962
rect 7986 11950 8016 11962
rect 8178 11950 8208 11962
rect 8370 11950 8400 11962
rect 8562 11950 8592 11962
rect 8754 11950 8784 11962
rect 9238 11950 9268 11962
rect 9430 11950 9460 11962
rect 9622 11950 9652 11962
rect 9814 11950 9844 11962
rect 10006 11950 10036 11962
rect 10198 11950 10228 11962
rect 10390 11950 10420 11962
rect 10582 11950 10612 11962
rect 11066 11950 11096 11962
rect 11258 11950 11288 11962
rect 11450 11950 11480 11962
rect 11642 11950 11672 11962
rect 11834 11950 11864 11962
rect 12026 11950 12056 11962
rect 12218 11950 12248 11962
rect 12410 11950 12440 11962
rect 12894 11950 12924 11962
rect 13086 11950 13116 11962
rect 13278 11950 13308 11962
rect 13470 11950 13500 11962
rect 13662 11950 13692 11962
rect 13854 11950 13884 11962
rect 14046 11950 14076 11962
rect 14238 11950 14268 11962
rect 14722 11950 14752 11962
rect 14914 11950 14944 11962
rect 15106 11950 15136 11962
rect 15298 11950 15328 11962
rect 15490 11950 15520 11962
rect 15682 11950 15712 11962
rect 15874 11950 15904 11962
rect 16066 11950 16096 11962
rect 16550 11950 16580 11962
rect 16742 11950 16772 11962
rect 16934 11950 16964 11962
rect 17126 11950 17156 11962
rect 17318 11950 17348 11962
rect 17510 11950 17540 11962
rect 17702 11950 17732 11962
rect 17894 11950 17924 11962
rect 18378 11950 18408 11962
rect 18570 11950 18600 11962
rect 18762 11950 18792 11962
rect 18954 11950 18984 11962
rect 19146 11950 19176 11962
rect 19338 11950 19368 11962
rect 19530 11950 19560 11962
rect 19722 11950 19752 11962
rect 20206 11950 20236 11962
rect 20398 11950 20428 11962
rect 20590 11950 20620 11962
rect 20782 11950 20812 11962
rect 20974 11950 21004 11962
rect 21166 11950 21196 11962
rect 21358 11950 21388 11962
rect 21550 11950 21580 11962
rect 194 11486 224 11498
rect 386 11486 416 11498
rect 578 11486 608 11498
rect 770 11486 800 11498
rect 962 11486 992 11498
rect 1154 11486 1184 11498
rect 1346 11486 1376 11498
rect 2022 11486 2052 11498
rect 2214 11486 2244 11498
rect 2406 11486 2436 11498
rect 2598 11486 2628 11498
rect 2790 11486 2820 11498
rect 2982 11486 3012 11498
rect 3174 11486 3204 11498
rect 3850 11486 3880 11498
rect 4042 11486 4072 11498
rect 4234 11486 4264 11498
rect 4426 11486 4456 11498
rect 4618 11486 4648 11498
rect 4810 11486 4840 11498
rect 5002 11486 5032 11498
rect 5678 11486 5708 11498
rect 5870 11486 5900 11498
rect 6062 11486 6092 11498
rect 6254 11486 6284 11498
rect 6446 11486 6476 11498
rect 6638 11486 6668 11498
rect 6830 11486 6860 11498
rect 7506 11486 7536 11498
rect 7698 11486 7728 11498
rect 7890 11486 7920 11498
rect 8082 11486 8112 11498
rect 8274 11486 8304 11498
rect 8466 11486 8496 11498
rect 8658 11486 8688 11498
rect 9334 11486 9364 11498
rect 9526 11486 9556 11498
rect 9718 11486 9748 11498
rect 9910 11486 9940 11498
rect 10102 11486 10132 11498
rect 10294 11486 10324 11498
rect 10486 11486 10516 11498
rect 11162 11486 11192 11498
rect 11354 11486 11384 11498
rect 11546 11486 11576 11498
rect 11738 11486 11768 11498
rect 11930 11486 11960 11498
rect 12122 11486 12152 11498
rect 12314 11486 12344 11498
rect 12990 11486 13020 11498
rect 13182 11486 13212 11498
rect 13374 11486 13404 11498
rect 13566 11486 13596 11498
rect 13758 11486 13788 11498
rect 13950 11486 13980 11498
rect 14142 11486 14172 11498
rect 14818 11486 14848 11498
rect 15010 11486 15040 11498
rect 15202 11486 15232 11498
rect 15394 11486 15424 11498
rect 15586 11486 15616 11498
rect 15778 11486 15808 11498
rect 15970 11486 16000 11498
rect 16646 11486 16676 11498
rect 16838 11486 16868 11498
rect 17030 11486 17060 11498
rect 17222 11486 17252 11498
rect 17414 11486 17444 11498
rect 17606 11486 17636 11498
rect 17798 11486 17828 11498
rect 18474 11486 18504 11498
rect 18666 11486 18696 11498
rect 18858 11486 18888 11498
rect 19050 11486 19080 11498
rect 19242 11486 19272 11498
rect 19434 11486 19464 11498
rect 19626 11486 19656 11498
rect 20302 11486 20332 11498
rect 20494 11486 20524 11498
rect 20686 11486 20716 11498
rect 20878 11486 20908 11498
rect 21070 11486 21100 11498
rect 21262 11486 21292 11498
rect 21454 11486 21484 11498
rect 0 11427 1490 11486
rect 1828 11427 3318 11486
rect 3656 11427 5146 11486
rect 5484 11427 6974 11486
rect 7312 11427 8802 11486
rect 9140 11427 10630 11486
rect 10968 11427 12458 11486
rect 12796 11427 14286 11486
rect 14624 11427 16114 11486
rect 16452 11427 17942 11486
rect 18280 11427 19770 11486
rect 20108 11427 21598 11486
rect 0 11248 1490 11307
rect 1828 11248 3318 11307
rect 3656 11248 5146 11307
rect 5484 11248 6974 11307
rect 7312 11248 8802 11307
rect 9140 11248 10630 11307
rect 10968 11248 12458 11307
rect 12796 11248 14286 11307
rect 14624 11248 16114 11307
rect 16452 11248 17942 11307
rect 18280 11248 19770 11307
rect 20108 11248 21598 11307
rect 98 11236 128 11248
rect 290 11236 320 11248
rect 482 11236 512 11248
rect 674 11236 704 11248
rect 866 11236 896 11248
rect 1058 11236 1088 11248
rect 1250 11236 1280 11248
rect 1442 11236 1472 11248
rect 1926 11236 1956 11248
rect 2118 11236 2148 11248
rect 2310 11236 2340 11248
rect 2502 11236 2532 11248
rect 2694 11236 2724 11248
rect 2886 11236 2916 11248
rect 3078 11236 3108 11248
rect 3270 11236 3300 11248
rect 3754 11236 3784 11248
rect 3946 11236 3976 11248
rect 4138 11236 4168 11248
rect 4330 11236 4360 11248
rect 4522 11236 4552 11248
rect 4714 11236 4744 11248
rect 4906 11236 4936 11248
rect 5098 11236 5128 11248
rect 5582 11236 5612 11248
rect 5774 11236 5804 11248
rect 5966 11236 5996 11248
rect 6158 11236 6188 11248
rect 6350 11236 6380 11248
rect 6542 11236 6572 11248
rect 6734 11236 6764 11248
rect 6926 11236 6956 11248
rect 7410 11236 7440 11248
rect 7602 11236 7632 11248
rect 7794 11236 7824 11248
rect 7986 11236 8016 11248
rect 8178 11236 8208 11248
rect 8370 11236 8400 11248
rect 8562 11236 8592 11248
rect 8754 11236 8784 11248
rect 9238 11236 9268 11248
rect 9430 11236 9460 11248
rect 9622 11236 9652 11248
rect 9814 11236 9844 11248
rect 10006 11236 10036 11248
rect 10198 11236 10228 11248
rect 10390 11236 10420 11248
rect 10582 11236 10612 11248
rect 11066 11236 11096 11248
rect 11258 11236 11288 11248
rect 11450 11236 11480 11248
rect 11642 11236 11672 11248
rect 11834 11236 11864 11248
rect 12026 11236 12056 11248
rect 12218 11236 12248 11248
rect 12410 11236 12440 11248
rect 12894 11236 12924 11248
rect 13086 11236 13116 11248
rect 13278 11236 13308 11248
rect 13470 11236 13500 11248
rect 13662 11236 13692 11248
rect 13854 11236 13884 11248
rect 14046 11236 14076 11248
rect 14238 11236 14268 11248
rect 14722 11236 14752 11248
rect 14914 11236 14944 11248
rect 15106 11236 15136 11248
rect 15298 11236 15328 11248
rect 15490 11236 15520 11248
rect 15682 11236 15712 11248
rect 15874 11236 15904 11248
rect 16066 11236 16096 11248
rect 16550 11236 16580 11248
rect 16742 11236 16772 11248
rect 16934 11236 16964 11248
rect 17126 11236 17156 11248
rect 17318 11236 17348 11248
rect 17510 11236 17540 11248
rect 17702 11236 17732 11248
rect 17894 11236 17924 11248
rect 18378 11236 18408 11248
rect 18570 11236 18600 11248
rect 18762 11236 18792 11248
rect 18954 11236 18984 11248
rect 19146 11236 19176 11248
rect 19338 11236 19368 11248
rect 19530 11236 19560 11248
rect 19722 11236 19752 11248
rect 20206 11236 20236 11248
rect 20398 11236 20428 11248
rect 20590 11236 20620 11248
rect 20782 11236 20812 11248
rect 20974 11236 21004 11248
rect 21166 11236 21196 11248
rect 21358 11236 21388 11248
rect 21550 11236 21580 11248
rect 194 10772 224 10784
rect 386 10772 416 10784
rect 578 10772 608 10784
rect 770 10772 800 10784
rect 962 10772 992 10784
rect 1154 10772 1184 10784
rect 1346 10772 1376 10784
rect 2022 10772 2052 10784
rect 2214 10772 2244 10784
rect 2406 10772 2436 10784
rect 2598 10772 2628 10784
rect 2790 10772 2820 10784
rect 2982 10772 3012 10784
rect 3174 10772 3204 10784
rect 3850 10772 3880 10784
rect 4042 10772 4072 10784
rect 4234 10772 4264 10784
rect 4426 10772 4456 10784
rect 4618 10772 4648 10784
rect 4810 10772 4840 10784
rect 5002 10772 5032 10784
rect 5678 10772 5708 10784
rect 5870 10772 5900 10784
rect 6062 10772 6092 10784
rect 6254 10772 6284 10784
rect 6446 10772 6476 10784
rect 6638 10772 6668 10784
rect 6830 10772 6860 10784
rect 7506 10772 7536 10784
rect 7698 10772 7728 10784
rect 7890 10772 7920 10784
rect 8082 10772 8112 10784
rect 8274 10772 8304 10784
rect 8466 10772 8496 10784
rect 8658 10772 8688 10784
rect 9334 10772 9364 10784
rect 9526 10772 9556 10784
rect 9718 10772 9748 10784
rect 9910 10772 9940 10784
rect 10102 10772 10132 10784
rect 10294 10772 10324 10784
rect 10486 10772 10516 10784
rect 11162 10772 11192 10784
rect 11354 10772 11384 10784
rect 11546 10772 11576 10784
rect 11738 10772 11768 10784
rect 11930 10772 11960 10784
rect 12122 10772 12152 10784
rect 12314 10772 12344 10784
rect 12990 10772 13020 10784
rect 13182 10772 13212 10784
rect 13374 10772 13404 10784
rect 13566 10772 13596 10784
rect 13758 10772 13788 10784
rect 13950 10772 13980 10784
rect 14142 10772 14172 10784
rect 14818 10772 14848 10784
rect 15010 10772 15040 10784
rect 15202 10772 15232 10784
rect 15394 10772 15424 10784
rect 15586 10772 15616 10784
rect 15778 10772 15808 10784
rect 15970 10772 16000 10784
rect 16646 10772 16676 10784
rect 16838 10772 16868 10784
rect 17030 10772 17060 10784
rect 17222 10772 17252 10784
rect 17414 10772 17444 10784
rect 17606 10772 17636 10784
rect 17798 10772 17828 10784
rect 18474 10772 18504 10784
rect 18666 10772 18696 10784
rect 18858 10772 18888 10784
rect 19050 10772 19080 10784
rect 19242 10772 19272 10784
rect 19434 10772 19464 10784
rect 19626 10772 19656 10784
rect 20302 10772 20332 10784
rect 20494 10772 20524 10784
rect 20686 10772 20716 10784
rect 20878 10772 20908 10784
rect 21070 10772 21100 10784
rect 21262 10772 21292 10784
rect 21454 10772 21484 10784
rect 0 10713 1490 10772
rect 1828 10713 3318 10772
rect 3656 10713 5146 10772
rect 5484 10713 6974 10772
rect 7312 10713 8802 10772
rect 9140 10713 10630 10772
rect 10968 10713 12458 10772
rect 12796 10713 14286 10772
rect 14624 10713 16114 10772
rect 16452 10713 17942 10772
rect 18280 10713 19770 10772
rect 20108 10713 21598 10772
rect 0 10534 1490 10593
rect 1828 10534 3318 10593
rect 3656 10534 5146 10593
rect 5484 10534 6974 10593
rect 7312 10534 8802 10593
rect 9140 10534 10630 10593
rect 10968 10534 12458 10593
rect 12796 10534 14286 10593
rect 14624 10534 16114 10593
rect 16452 10534 17942 10593
rect 18280 10534 19770 10593
rect 20108 10534 21598 10593
rect 98 10522 128 10534
rect 290 10522 320 10534
rect 482 10522 512 10534
rect 674 10522 704 10534
rect 866 10522 896 10534
rect 1058 10522 1088 10534
rect 1250 10522 1280 10534
rect 1442 10522 1472 10534
rect 1926 10522 1956 10534
rect 2118 10522 2148 10534
rect 2310 10522 2340 10534
rect 2502 10522 2532 10534
rect 2694 10522 2724 10534
rect 2886 10522 2916 10534
rect 3078 10522 3108 10534
rect 3270 10522 3300 10534
rect 3754 10522 3784 10534
rect 3946 10522 3976 10534
rect 4138 10522 4168 10534
rect 4330 10522 4360 10534
rect 4522 10522 4552 10534
rect 4714 10522 4744 10534
rect 4906 10522 4936 10534
rect 5098 10522 5128 10534
rect 5582 10522 5612 10534
rect 5774 10522 5804 10534
rect 5966 10522 5996 10534
rect 6158 10522 6188 10534
rect 6350 10522 6380 10534
rect 6542 10522 6572 10534
rect 6734 10522 6764 10534
rect 6926 10522 6956 10534
rect 7410 10522 7440 10534
rect 7602 10522 7632 10534
rect 7794 10522 7824 10534
rect 7986 10522 8016 10534
rect 8178 10522 8208 10534
rect 8370 10522 8400 10534
rect 8562 10522 8592 10534
rect 8754 10522 8784 10534
rect 9238 10522 9268 10534
rect 9430 10522 9460 10534
rect 9622 10522 9652 10534
rect 9814 10522 9844 10534
rect 10006 10522 10036 10534
rect 10198 10522 10228 10534
rect 10390 10522 10420 10534
rect 10582 10522 10612 10534
rect 11066 10522 11096 10534
rect 11258 10522 11288 10534
rect 11450 10522 11480 10534
rect 11642 10522 11672 10534
rect 11834 10522 11864 10534
rect 12026 10522 12056 10534
rect 12218 10522 12248 10534
rect 12410 10522 12440 10534
rect 12894 10522 12924 10534
rect 13086 10522 13116 10534
rect 13278 10522 13308 10534
rect 13470 10522 13500 10534
rect 13662 10522 13692 10534
rect 13854 10522 13884 10534
rect 14046 10522 14076 10534
rect 14238 10522 14268 10534
rect 14722 10522 14752 10534
rect 14914 10522 14944 10534
rect 15106 10522 15136 10534
rect 15298 10522 15328 10534
rect 15490 10522 15520 10534
rect 15682 10522 15712 10534
rect 15874 10522 15904 10534
rect 16066 10522 16096 10534
rect 16550 10522 16580 10534
rect 16742 10522 16772 10534
rect 16934 10522 16964 10534
rect 17126 10522 17156 10534
rect 17318 10522 17348 10534
rect 17510 10522 17540 10534
rect 17702 10522 17732 10534
rect 17894 10522 17924 10534
rect 18378 10522 18408 10534
rect 18570 10522 18600 10534
rect 18762 10522 18792 10534
rect 18954 10522 18984 10534
rect 19146 10522 19176 10534
rect 19338 10522 19368 10534
rect 19530 10522 19560 10534
rect 19722 10522 19752 10534
rect 20206 10522 20236 10534
rect 20398 10522 20428 10534
rect 20590 10522 20620 10534
rect 20782 10522 20812 10534
rect 20974 10522 21004 10534
rect 21166 10522 21196 10534
rect 21358 10522 21388 10534
rect 21550 10522 21580 10534
rect 194 10058 224 10070
rect 386 10058 416 10070
rect 578 10058 608 10070
rect 770 10058 800 10070
rect 962 10058 992 10070
rect 1154 10058 1184 10070
rect 1346 10058 1376 10070
rect 2022 10058 2052 10070
rect 2214 10058 2244 10070
rect 2406 10058 2436 10070
rect 2598 10058 2628 10070
rect 2790 10058 2820 10070
rect 2982 10058 3012 10070
rect 3174 10058 3204 10070
rect 3850 10058 3880 10070
rect 4042 10058 4072 10070
rect 4234 10058 4264 10070
rect 4426 10058 4456 10070
rect 4618 10058 4648 10070
rect 4810 10058 4840 10070
rect 5002 10058 5032 10070
rect 5678 10058 5708 10070
rect 5870 10058 5900 10070
rect 6062 10058 6092 10070
rect 6254 10058 6284 10070
rect 6446 10058 6476 10070
rect 6638 10058 6668 10070
rect 6830 10058 6860 10070
rect 7506 10058 7536 10070
rect 7698 10058 7728 10070
rect 7890 10058 7920 10070
rect 8082 10058 8112 10070
rect 8274 10058 8304 10070
rect 8466 10058 8496 10070
rect 8658 10058 8688 10070
rect 9334 10058 9364 10070
rect 9526 10058 9556 10070
rect 9718 10058 9748 10070
rect 9910 10058 9940 10070
rect 10102 10058 10132 10070
rect 10294 10058 10324 10070
rect 10486 10058 10516 10070
rect 11162 10058 11192 10070
rect 11354 10058 11384 10070
rect 11546 10058 11576 10070
rect 11738 10058 11768 10070
rect 11930 10058 11960 10070
rect 12122 10058 12152 10070
rect 12314 10058 12344 10070
rect 12990 10058 13020 10070
rect 13182 10058 13212 10070
rect 13374 10058 13404 10070
rect 13566 10058 13596 10070
rect 13758 10058 13788 10070
rect 13950 10058 13980 10070
rect 14142 10058 14172 10070
rect 14818 10058 14848 10070
rect 15010 10058 15040 10070
rect 15202 10058 15232 10070
rect 15394 10058 15424 10070
rect 15586 10058 15616 10070
rect 15778 10058 15808 10070
rect 15970 10058 16000 10070
rect 16646 10058 16676 10070
rect 16838 10058 16868 10070
rect 17030 10058 17060 10070
rect 17222 10058 17252 10070
rect 17414 10058 17444 10070
rect 17606 10058 17636 10070
rect 17798 10058 17828 10070
rect 18474 10058 18504 10070
rect 18666 10058 18696 10070
rect 18858 10058 18888 10070
rect 19050 10058 19080 10070
rect 19242 10058 19272 10070
rect 19434 10058 19464 10070
rect 19626 10058 19656 10070
rect 20302 10058 20332 10070
rect 20494 10058 20524 10070
rect 20686 10058 20716 10070
rect 20878 10058 20908 10070
rect 21070 10058 21100 10070
rect 21262 10058 21292 10070
rect 21454 10058 21484 10070
rect 0 9999 1490 10058
rect 1828 9999 3318 10058
rect 3656 9999 5146 10058
rect 5484 9999 6974 10058
rect 7312 9999 8802 10058
rect 9140 9999 10630 10058
rect 10968 9999 12458 10058
rect 12796 9999 14286 10058
rect 14624 9999 16114 10058
rect 16452 9999 17942 10058
rect 18280 9999 19770 10058
rect 20108 9999 21598 10058
rect 0 9820 1490 9879
rect 1828 9820 3318 9879
rect 3656 9820 5146 9879
rect 5484 9820 6974 9879
rect 7312 9820 8802 9879
rect 9140 9820 10630 9879
rect 10968 9820 12458 9879
rect 12796 9820 14286 9879
rect 14624 9820 16114 9879
rect 16452 9820 17942 9879
rect 18280 9820 19770 9879
rect 20108 9820 21598 9879
rect 98 9808 128 9820
rect 290 9808 320 9820
rect 482 9808 512 9820
rect 674 9808 704 9820
rect 866 9808 896 9820
rect 1058 9808 1088 9820
rect 1250 9808 1280 9820
rect 1442 9808 1472 9820
rect 1926 9808 1956 9820
rect 2118 9808 2148 9820
rect 2310 9808 2340 9820
rect 2502 9808 2532 9820
rect 2694 9808 2724 9820
rect 2886 9808 2916 9820
rect 3078 9808 3108 9820
rect 3270 9808 3300 9820
rect 3754 9808 3784 9820
rect 3946 9808 3976 9820
rect 4138 9808 4168 9820
rect 4330 9808 4360 9820
rect 4522 9808 4552 9820
rect 4714 9808 4744 9820
rect 4906 9808 4936 9820
rect 5098 9808 5128 9820
rect 5582 9808 5612 9820
rect 5774 9808 5804 9820
rect 5966 9808 5996 9820
rect 6158 9808 6188 9820
rect 6350 9808 6380 9820
rect 6542 9808 6572 9820
rect 6734 9808 6764 9820
rect 6926 9808 6956 9820
rect 7410 9808 7440 9820
rect 7602 9808 7632 9820
rect 7794 9808 7824 9820
rect 7986 9808 8016 9820
rect 8178 9808 8208 9820
rect 8370 9808 8400 9820
rect 8562 9808 8592 9820
rect 8754 9808 8784 9820
rect 9238 9808 9268 9820
rect 9430 9808 9460 9820
rect 9622 9808 9652 9820
rect 9814 9808 9844 9820
rect 10006 9808 10036 9820
rect 10198 9808 10228 9820
rect 10390 9808 10420 9820
rect 10582 9808 10612 9820
rect 11066 9808 11096 9820
rect 11258 9808 11288 9820
rect 11450 9808 11480 9820
rect 11642 9808 11672 9820
rect 11834 9808 11864 9820
rect 12026 9808 12056 9820
rect 12218 9808 12248 9820
rect 12410 9808 12440 9820
rect 12894 9808 12924 9820
rect 13086 9808 13116 9820
rect 13278 9808 13308 9820
rect 13470 9808 13500 9820
rect 13662 9808 13692 9820
rect 13854 9808 13884 9820
rect 14046 9808 14076 9820
rect 14238 9808 14268 9820
rect 14722 9808 14752 9820
rect 14914 9808 14944 9820
rect 15106 9808 15136 9820
rect 15298 9808 15328 9820
rect 15490 9808 15520 9820
rect 15682 9808 15712 9820
rect 15874 9808 15904 9820
rect 16066 9808 16096 9820
rect 16550 9808 16580 9820
rect 16742 9808 16772 9820
rect 16934 9808 16964 9820
rect 17126 9808 17156 9820
rect 17318 9808 17348 9820
rect 17510 9808 17540 9820
rect 17702 9808 17732 9820
rect 17894 9808 17924 9820
rect 18378 9808 18408 9820
rect 18570 9808 18600 9820
rect 18762 9808 18792 9820
rect 18954 9808 18984 9820
rect 19146 9808 19176 9820
rect 19338 9808 19368 9820
rect 19530 9808 19560 9820
rect 19722 9808 19752 9820
rect 20206 9808 20236 9820
rect 20398 9808 20428 9820
rect 20590 9808 20620 9820
rect 20782 9808 20812 9820
rect 20974 9808 21004 9820
rect 21166 9808 21196 9820
rect 21358 9808 21388 9820
rect 21550 9808 21580 9820
rect 194 9344 224 9356
rect 386 9344 416 9356
rect 578 9344 608 9356
rect 770 9344 800 9356
rect 962 9344 992 9356
rect 1154 9344 1184 9356
rect 1346 9344 1376 9356
rect 2022 9344 2052 9356
rect 2214 9344 2244 9356
rect 2406 9344 2436 9356
rect 2598 9344 2628 9356
rect 2790 9344 2820 9356
rect 2982 9344 3012 9356
rect 3174 9344 3204 9356
rect 3850 9344 3880 9356
rect 4042 9344 4072 9356
rect 4234 9344 4264 9356
rect 4426 9344 4456 9356
rect 4618 9344 4648 9356
rect 4810 9344 4840 9356
rect 5002 9344 5032 9356
rect 5678 9344 5708 9356
rect 5870 9344 5900 9356
rect 6062 9344 6092 9356
rect 6254 9344 6284 9356
rect 6446 9344 6476 9356
rect 6638 9344 6668 9356
rect 6830 9344 6860 9356
rect 7506 9344 7536 9356
rect 7698 9344 7728 9356
rect 7890 9344 7920 9356
rect 8082 9344 8112 9356
rect 8274 9344 8304 9356
rect 8466 9344 8496 9356
rect 8658 9344 8688 9356
rect 9334 9344 9364 9356
rect 9526 9344 9556 9356
rect 9718 9344 9748 9356
rect 9910 9344 9940 9356
rect 10102 9344 10132 9356
rect 10294 9344 10324 9356
rect 10486 9344 10516 9356
rect 11162 9344 11192 9356
rect 11354 9344 11384 9356
rect 11546 9344 11576 9356
rect 11738 9344 11768 9356
rect 11930 9344 11960 9356
rect 12122 9344 12152 9356
rect 12314 9344 12344 9356
rect 12990 9344 13020 9356
rect 13182 9344 13212 9356
rect 13374 9344 13404 9356
rect 13566 9344 13596 9356
rect 13758 9344 13788 9356
rect 13950 9344 13980 9356
rect 14142 9344 14172 9356
rect 14818 9344 14848 9356
rect 15010 9344 15040 9356
rect 15202 9344 15232 9356
rect 15394 9344 15424 9356
rect 15586 9344 15616 9356
rect 15778 9344 15808 9356
rect 15970 9344 16000 9356
rect 16646 9344 16676 9356
rect 16838 9344 16868 9356
rect 17030 9344 17060 9356
rect 17222 9344 17252 9356
rect 17414 9344 17444 9356
rect 17606 9344 17636 9356
rect 17798 9344 17828 9356
rect 18474 9344 18504 9356
rect 18666 9344 18696 9356
rect 18858 9344 18888 9356
rect 19050 9344 19080 9356
rect 19242 9344 19272 9356
rect 19434 9344 19464 9356
rect 19626 9344 19656 9356
rect 20302 9344 20332 9356
rect 20494 9344 20524 9356
rect 20686 9344 20716 9356
rect 20878 9344 20908 9356
rect 21070 9344 21100 9356
rect 21262 9344 21292 9356
rect 21454 9344 21484 9356
rect 0 9285 1490 9344
rect 1828 9285 3318 9344
rect 3656 9285 5146 9344
rect 5484 9285 6974 9344
rect 7312 9285 8802 9344
rect 9140 9285 10630 9344
rect 10968 9285 12458 9344
rect 12796 9285 14286 9344
rect 14624 9285 16114 9344
rect 16452 9285 17942 9344
rect 18280 9285 19770 9344
rect 20108 9285 21598 9344
rect 0 9106 1490 9165
rect 1828 9106 3318 9165
rect 3656 9106 5146 9165
rect 5484 9106 6974 9165
rect 7312 9106 8802 9165
rect 9140 9106 10630 9165
rect 10968 9106 12458 9165
rect 12796 9106 14286 9165
rect 14624 9106 16114 9165
rect 16452 9106 17942 9165
rect 18280 9106 19770 9165
rect 20108 9106 21598 9165
rect 98 9094 128 9106
rect 290 9094 320 9106
rect 482 9094 512 9106
rect 674 9094 704 9106
rect 866 9094 896 9106
rect 1058 9094 1088 9106
rect 1250 9094 1280 9106
rect 1442 9094 1472 9106
rect 1926 9094 1956 9106
rect 2118 9094 2148 9106
rect 2310 9094 2340 9106
rect 2502 9094 2532 9106
rect 2694 9094 2724 9106
rect 2886 9094 2916 9106
rect 3078 9094 3108 9106
rect 3270 9094 3300 9106
rect 3754 9094 3784 9106
rect 3946 9094 3976 9106
rect 4138 9094 4168 9106
rect 4330 9094 4360 9106
rect 4522 9094 4552 9106
rect 4714 9094 4744 9106
rect 4906 9094 4936 9106
rect 5098 9094 5128 9106
rect 5582 9094 5612 9106
rect 5774 9094 5804 9106
rect 5966 9094 5996 9106
rect 6158 9094 6188 9106
rect 6350 9094 6380 9106
rect 6542 9094 6572 9106
rect 6734 9094 6764 9106
rect 6926 9094 6956 9106
rect 7410 9094 7440 9106
rect 7602 9094 7632 9106
rect 7794 9094 7824 9106
rect 7986 9094 8016 9106
rect 8178 9094 8208 9106
rect 8370 9094 8400 9106
rect 8562 9094 8592 9106
rect 8754 9094 8784 9106
rect 9238 9094 9268 9106
rect 9430 9094 9460 9106
rect 9622 9094 9652 9106
rect 9814 9094 9844 9106
rect 10006 9094 10036 9106
rect 10198 9094 10228 9106
rect 10390 9094 10420 9106
rect 10582 9094 10612 9106
rect 11066 9094 11096 9106
rect 11258 9094 11288 9106
rect 11450 9094 11480 9106
rect 11642 9094 11672 9106
rect 11834 9094 11864 9106
rect 12026 9094 12056 9106
rect 12218 9094 12248 9106
rect 12410 9094 12440 9106
rect 12894 9094 12924 9106
rect 13086 9094 13116 9106
rect 13278 9094 13308 9106
rect 13470 9094 13500 9106
rect 13662 9094 13692 9106
rect 13854 9094 13884 9106
rect 14046 9094 14076 9106
rect 14238 9094 14268 9106
rect 14722 9094 14752 9106
rect 14914 9094 14944 9106
rect 15106 9094 15136 9106
rect 15298 9094 15328 9106
rect 15490 9094 15520 9106
rect 15682 9094 15712 9106
rect 15874 9094 15904 9106
rect 16066 9094 16096 9106
rect 16550 9094 16580 9106
rect 16742 9094 16772 9106
rect 16934 9094 16964 9106
rect 17126 9094 17156 9106
rect 17318 9094 17348 9106
rect 17510 9094 17540 9106
rect 17702 9094 17732 9106
rect 17894 9094 17924 9106
rect 18378 9094 18408 9106
rect 18570 9094 18600 9106
rect 18762 9094 18792 9106
rect 18954 9094 18984 9106
rect 19146 9094 19176 9106
rect 19338 9094 19368 9106
rect 19530 9094 19560 9106
rect 19722 9094 19752 9106
rect 20206 9094 20236 9106
rect 20398 9094 20428 9106
rect 20590 9094 20620 9106
rect 20782 9094 20812 9106
rect 20974 9094 21004 9106
rect 21166 9094 21196 9106
rect 21358 9094 21388 9106
rect 21550 9094 21580 9106
rect 194 8630 224 8642
rect 386 8630 416 8642
rect 578 8630 608 8642
rect 770 8630 800 8642
rect 962 8630 992 8642
rect 1154 8630 1184 8642
rect 1346 8630 1376 8642
rect 2022 8630 2052 8642
rect 2214 8630 2244 8642
rect 2406 8630 2436 8642
rect 2598 8630 2628 8642
rect 2790 8630 2820 8642
rect 2982 8630 3012 8642
rect 3174 8630 3204 8642
rect 3850 8630 3880 8642
rect 4042 8630 4072 8642
rect 4234 8630 4264 8642
rect 4426 8630 4456 8642
rect 4618 8630 4648 8642
rect 4810 8630 4840 8642
rect 5002 8630 5032 8642
rect 5678 8630 5708 8642
rect 5870 8630 5900 8642
rect 6062 8630 6092 8642
rect 6254 8630 6284 8642
rect 6446 8630 6476 8642
rect 6638 8630 6668 8642
rect 6830 8630 6860 8642
rect 7506 8630 7536 8642
rect 7698 8630 7728 8642
rect 7890 8630 7920 8642
rect 8082 8630 8112 8642
rect 8274 8630 8304 8642
rect 8466 8630 8496 8642
rect 8658 8630 8688 8642
rect 9334 8630 9364 8642
rect 9526 8630 9556 8642
rect 9718 8630 9748 8642
rect 9910 8630 9940 8642
rect 10102 8630 10132 8642
rect 10294 8630 10324 8642
rect 10486 8630 10516 8642
rect 11162 8630 11192 8642
rect 11354 8630 11384 8642
rect 11546 8630 11576 8642
rect 11738 8630 11768 8642
rect 11930 8630 11960 8642
rect 12122 8630 12152 8642
rect 12314 8630 12344 8642
rect 12990 8630 13020 8642
rect 13182 8630 13212 8642
rect 13374 8630 13404 8642
rect 13566 8630 13596 8642
rect 13758 8630 13788 8642
rect 13950 8630 13980 8642
rect 14142 8630 14172 8642
rect 14818 8630 14848 8642
rect 15010 8630 15040 8642
rect 15202 8630 15232 8642
rect 15394 8630 15424 8642
rect 15586 8630 15616 8642
rect 15778 8630 15808 8642
rect 15970 8630 16000 8642
rect 16646 8630 16676 8642
rect 16838 8630 16868 8642
rect 17030 8630 17060 8642
rect 17222 8630 17252 8642
rect 17414 8630 17444 8642
rect 17606 8630 17636 8642
rect 17798 8630 17828 8642
rect 18474 8630 18504 8642
rect 18666 8630 18696 8642
rect 18858 8630 18888 8642
rect 19050 8630 19080 8642
rect 19242 8630 19272 8642
rect 19434 8630 19464 8642
rect 19626 8630 19656 8642
rect 20302 8630 20332 8642
rect 20494 8630 20524 8642
rect 20686 8630 20716 8642
rect 20878 8630 20908 8642
rect 21070 8630 21100 8642
rect 21262 8630 21292 8642
rect 21454 8630 21484 8642
rect 0 8571 1490 8630
rect 1828 8571 3318 8630
rect 3656 8571 5146 8630
rect 5484 8571 6974 8630
rect 7312 8571 8802 8630
rect 9140 8571 10630 8630
rect 10968 8571 12458 8630
rect 12796 8571 14286 8630
rect 14624 8571 16114 8630
rect 16452 8571 17942 8630
rect 18280 8571 19770 8630
rect 20108 8571 21598 8630
rect 0 8392 1490 8451
rect 1828 8392 3318 8451
rect 3656 8392 5146 8451
rect 5484 8392 6974 8451
rect 7312 8392 8802 8451
rect 9140 8392 10630 8451
rect 10968 8392 12458 8451
rect 12796 8392 14286 8451
rect 14624 8392 16114 8451
rect 16452 8392 17942 8451
rect 18280 8392 19770 8451
rect 20108 8392 21598 8451
rect 98 8380 128 8392
rect 290 8380 320 8392
rect 482 8380 512 8392
rect 674 8380 704 8392
rect 866 8380 896 8392
rect 1058 8380 1088 8392
rect 1250 8380 1280 8392
rect 1442 8380 1472 8392
rect 1926 8380 1956 8392
rect 2118 8380 2148 8392
rect 2310 8380 2340 8392
rect 2502 8380 2532 8392
rect 2694 8380 2724 8392
rect 2886 8380 2916 8392
rect 3078 8380 3108 8392
rect 3270 8380 3300 8392
rect 3754 8380 3784 8392
rect 3946 8380 3976 8392
rect 4138 8380 4168 8392
rect 4330 8380 4360 8392
rect 4522 8380 4552 8392
rect 4714 8380 4744 8392
rect 4906 8380 4936 8392
rect 5098 8380 5128 8392
rect 5582 8380 5612 8392
rect 5774 8380 5804 8392
rect 5966 8380 5996 8392
rect 6158 8380 6188 8392
rect 6350 8380 6380 8392
rect 6542 8380 6572 8392
rect 6734 8380 6764 8392
rect 6926 8380 6956 8392
rect 7410 8380 7440 8392
rect 7602 8380 7632 8392
rect 7794 8380 7824 8392
rect 7986 8380 8016 8392
rect 8178 8380 8208 8392
rect 8370 8380 8400 8392
rect 8562 8380 8592 8392
rect 8754 8380 8784 8392
rect 9238 8380 9268 8392
rect 9430 8380 9460 8392
rect 9622 8380 9652 8392
rect 9814 8380 9844 8392
rect 10006 8380 10036 8392
rect 10198 8380 10228 8392
rect 10390 8380 10420 8392
rect 10582 8380 10612 8392
rect 11066 8380 11096 8392
rect 11258 8380 11288 8392
rect 11450 8380 11480 8392
rect 11642 8380 11672 8392
rect 11834 8380 11864 8392
rect 12026 8380 12056 8392
rect 12218 8380 12248 8392
rect 12410 8380 12440 8392
rect 12894 8380 12924 8392
rect 13086 8380 13116 8392
rect 13278 8380 13308 8392
rect 13470 8380 13500 8392
rect 13662 8380 13692 8392
rect 13854 8380 13884 8392
rect 14046 8380 14076 8392
rect 14238 8380 14268 8392
rect 14722 8380 14752 8392
rect 14914 8380 14944 8392
rect 15106 8380 15136 8392
rect 15298 8380 15328 8392
rect 15490 8380 15520 8392
rect 15682 8380 15712 8392
rect 15874 8380 15904 8392
rect 16066 8380 16096 8392
rect 16550 8380 16580 8392
rect 16742 8380 16772 8392
rect 16934 8380 16964 8392
rect 17126 8380 17156 8392
rect 17318 8380 17348 8392
rect 17510 8380 17540 8392
rect 17702 8380 17732 8392
rect 17894 8380 17924 8392
rect 18378 8380 18408 8392
rect 18570 8380 18600 8392
rect 18762 8380 18792 8392
rect 18954 8380 18984 8392
rect 19146 8380 19176 8392
rect 19338 8380 19368 8392
rect 19530 8380 19560 8392
rect 19722 8380 19752 8392
rect 20206 8380 20236 8392
rect 20398 8380 20428 8392
rect 20590 8380 20620 8392
rect 20782 8380 20812 8392
rect 20974 8380 21004 8392
rect 21166 8380 21196 8392
rect 21358 8380 21388 8392
rect 21550 8380 21580 8392
rect 194 7916 224 7928
rect 386 7916 416 7928
rect 578 7916 608 7928
rect 770 7916 800 7928
rect 962 7916 992 7928
rect 1154 7916 1184 7928
rect 1346 7916 1376 7928
rect 2022 7916 2052 7928
rect 2214 7916 2244 7928
rect 2406 7916 2436 7928
rect 2598 7916 2628 7928
rect 2790 7916 2820 7928
rect 2982 7916 3012 7928
rect 3174 7916 3204 7928
rect 3850 7916 3880 7928
rect 4042 7916 4072 7928
rect 4234 7916 4264 7928
rect 4426 7916 4456 7928
rect 4618 7916 4648 7928
rect 4810 7916 4840 7928
rect 5002 7916 5032 7928
rect 5678 7916 5708 7928
rect 5870 7916 5900 7928
rect 6062 7916 6092 7928
rect 6254 7916 6284 7928
rect 6446 7916 6476 7928
rect 6638 7916 6668 7928
rect 6830 7916 6860 7928
rect 7506 7916 7536 7928
rect 7698 7916 7728 7928
rect 7890 7916 7920 7928
rect 8082 7916 8112 7928
rect 8274 7916 8304 7928
rect 8466 7916 8496 7928
rect 8658 7916 8688 7928
rect 9334 7916 9364 7928
rect 9526 7916 9556 7928
rect 9718 7916 9748 7928
rect 9910 7916 9940 7928
rect 10102 7916 10132 7928
rect 10294 7916 10324 7928
rect 10486 7916 10516 7928
rect 11162 7916 11192 7928
rect 11354 7916 11384 7928
rect 11546 7916 11576 7928
rect 11738 7916 11768 7928
rect 11930 7916 11960 7928
rect 12122 7916 12152 7928
rect 12314 7916 12344 7928
rect 12990 7916 13020 7928
rect 13182 7916 13212 7928
rect 13374 7916 13404 7928
rect 13566 7916 13596 7928
rect 13758 7916 13788 7928
rect 13950 7916 13980 7928
rect 14142 7916 14172 7928
rect 14818 7916 14848 7928
rect 15010 7916 15040 7928
rect 15202 7916 15232 7928
rect 15394 7916 15424 7928
rect 15586 7916 15616 7928
rect 15778 7916 15808 7928
rect 15970 7916 16000 7928
rect 16646 7916 16676 7928
rect 16838 7916 16868 7928
rect 17030 7916 17060 7928
rect 17222 7916 17252 7928
rect 17414 7916 17444 7928
rect 17606 7916 17636 7928
rect 17798 7916 17828 7928
rect 18474 7916 18504 7928
rect 18666 7916 18696 7928
rect 18858 7916 18888 7928
rect 19050 7916 19080 7928
rect 19242 7916 19272 7928
rect 19434 7916 19464 7928
rect 19626 7916 19656 7928
rect 20302 7916 20332 7928
rect 20494 7916 20524 7928
rect 20686 7916 20716 7928
rect 20878 7916 20908 7928
rect 21070 7916 21100 7928
rect 21262 7916 21292 7928
rect 21454 7916 21484 7928
rect 0 7857 1490 7916
rect 1828 7857 3318 7916
rect 3656 7857 5146 7916
rect 5484 7857 6974 7916
rect 7312 7857 8802 7916
rect 9140 7857 10630 7916
rect 10968 7857 12458 7916
rect 12796 7857 14286 7916
rect 14624 7857 16114 7916
rect 16452 7857 17942 7916
rect 18280 7857 19770 7916
rect 20108 7857 21598 7916
rect 0 7678 1490 7737
rect 1828 7678 3318 7737
rect 3656 7678 5146 7737
rect 5484 7678 6974 7737
rect 7312 7678 8802 7737
rect 9140 7678 10630 7737
rect 10968 7678 12458 7737
rect 12796 7678 14286 7737
rect 14624 7678 16114 7737
rect 16452 7678 17942 7737
rect 18280 7678 19770 7737
rect 20108 7678 21598 7737
rect 98 7666 128 7678
rect 290 7666 320 7678
rect 482 7666 512 7678
rect 674 7666 704 7678
rect 866 7666 896 7678
rect 1058 7666 1088 7678
rect 1250 7666 1280 7678
rect 1442 7666 1472 7678
rect 1926 7666 1956 7678
rect 2118 7666 2148 7678
rect 2310 7666 2340 7678
rect 2502 7666 2532 7678
rect 2694 7666 2724 7678
rect 2886 7666 2916 7678
rect 3078 7666 3108 7678
rect 3270 7666 3300 7678
rect 3754 7666 3784 7678
rect 3946 7666 3976 7678
rect 4138 7666 4168 7678
rect 4330 7666 4360 7678
rect 4522 7666 4552 7678
rect 4714 7666 4744 7678
rect 4906 7666 4936 7678
rect 5098 7666 5128 7678
rect 5582 7666 5612 7678
rect 5774 7666 5804 7678
rect 5966 7666 5996 7678
rect 6158 7666 6188 7678
rect 6350 7666 6380 7678
rect 6542 7666 6572 7678
rect 6734 7666 6764 7678
rect 6926 7666 6956 7678
rect 7410 7666 7440 7678
rect 7602 7666 7632 7678
rect 7794 7666 7824 7678
rect 7986 7666 8016 7678
rect 8178 7666 8208 7678
rect 8370 7666 8400 7678
rect 8562 7666 8592 7678
rect 8754 7666 8784 7678
rect 9238 7666 9268 7678
rect 9430 7666 9460 7678
rect 9622 7666 9652 7678
rect 9814 7666 9844 7678
rect 10006 7666 10036 7678
rect 10198 7666 10228 7678
rect 10390 7666 10420 7678
rect 10582 7666 10612 7678
rect 11066 7666 11096 7678
rect 11258 7666 11288 7678
rect 11450 7666 11480 7678
rect 11642 7666 11672 7678
rect 11834 7666 11864 7678
rect 12026 7666 12056 7678
rect 12218 7666 12248 7678
rect 12410 7666 12440 7678
rect 12894 7666 12924 7678
rect 13086 7666 13116 7678
rect 13278 7666 13308 7678
rect 13470 7666 13500 7678
rect 13662 7666 13692 7678
rect 13854 7666 13884 7678
rect 14046 7666 14076 7678
rect 14238 7666 14268 7678
rect 14722 7666 14752 7678
rect 14914 7666 14944 7678
rect 15106 7666 15136 7678
rect 15298 7666 15328 7678
rect 15490 7666 15520 7678
rect 15682 7666 15712 7678
rect 15874 7666 15904 7678
rect 16066 7666 16096 7678
rect 16550 7666 16580 7678
rect 16742 7666 16772 7678
rect 16934 7666 16964 7678
rect 17126 7666 17156 7678
rect 17318 7666 17348 7678
rect 17510 7666 17540 7678
rect 17702 7666 17732 7678
rect 17894 7666 17924 7678
rect 18378 7666 18408 7678
rect 18570 7666 18600 7678
rect 18762 7666 18792 7678
rect 18954 7666 18984 7678
rect 19146 7666 19176 7678
rect 19338 7666 19368 7678
rect 19530 7666 19560 7678
rect 19722 7666 19752 7678
rect 20206 7666 20236 7678
rect 20398 7666 20428 7678
rect 20590 7666 20620 7678
rect 20782 7666 20812 7678
rect 20974 7666 21004 7678
rect 21166 7666 21196 7678
rect 21358 7666 21388 7678
rect 21550 7666 21580 7678
rect 194 7202 224 7214
rect 386 7202 416 7214
rect 578 7202 608 7214
rect 770 7202 800 7214
rect 962 7202 992 7214
rect 1154 7202 1184 7214
rect 1346 7202 1376 7214
rect 2022 7202 2052 7214
rect 2214 7202 2244 7214
rect 2406 7202 2436 7214
rect 2598 7202 2628 7214
rect 2790 7202 2820 7214
rect 2982 7202 3012 7214
rect 3174 7202 3204 7214
rect 3850 7202 3880 7214
rect 4042 7202 4072 7214
rect 4234 7202 4264 7214
rect 4426 7202 4456 7214
rect 4618 7202 4648 7214
rect 4810 7202 4840 7214
rect 5002 7202 5032 7214
rect 5678 7202 5708 7214
rect 5870 7202 5900 7214
rect 6062 7202 6092 7214
rect 6254 7202 6284 7214
rect 6446 7202 6476 7214
rect 6638 7202 6668 7214
rect 6830 7202 6860 7214
rect 7506 7202 7536 7214
rect 7698 7202 7728 7214
rect 7890 7202 7920 7214
rect 8082 7202 8112 7214
rect 8274 7202 8304 7214
rect 8466 7202 8496 7214
rect 8658 7202 8688 7214
rect 9334 7202 9364 7214
rect 9526 7202 9556 7214
rect 9718 7202 9748 7214
rect 9910 7202 9940 7214
rect 10102 7202 10132 7214
rect 10294 7202 10324 7214
rect 10486 7202 10516 7214
rect 11162 7202 11192 7214
rect 11354 7202 11384 7214
rect 11546 7202 11576 7214
rect 11738 7202 11768 7214
rect 11930 7202 11960 7214
rect 12122 7202 12152 7214
rect 12314 7202 12344 7214
rect 12990 7202 13020 7214
rect 13182 7202 13212 7214
rect 13374 7202 13404 7214
rect 13566 7202 13596 7214
rect 13758 7202 13788 7214
rect 13950 7202 13980 7214
rect 14142 7202 14172 7214
rect 14818 7202 14848 7214
rect 15010 7202 15040 7214
rect 15202 7202 15232 7214
rect 15394 7202 15424 7214
rect 15586 7202 15616 7214
rect 15778 7202 15808 7214
rect 15970 7202 16000 7214
rect 16646 7202 16676 7214
rect 16838 7202 16868 7214
rect 17030 7202 17060 7214
rect 17222 7202 17252 7214
rect 17414 7202 17444 7214
rect 17606 7202 17636 7214
rect 17798 7202 17828 7214
rect 18474 7202 18504 7214
rect 18666 7202 18696 7214
rect 18858 7202 18888 7214
rect 19050 7202 19080 7214
rect 19242 7202 19272 7214
rect 19434 7202 19464 7214
rect 19626 7202 19656 7214
rect 20302 7202 20332 7214
rect 20494 7202 20524 7214
rect 20686 7202 20716 7214
rect 20878 7202 20908 7214
rect 21070 7202 21100 7214
rect 21262 7202 21292 7214
rect 21454 7202 21484 7214
rect 0 7143 1490 7202
rect 1828 7143 3318 7202
rect 3656 7143 5146 7202
rect 5484 7143 6974 7202
rect 7312 7143 8802 7202
rect 9140 7143 10630 7202
rect 10968 7143 12458 7202
rect 12796 7143 14286 7202
rect 14624 7143 16114 7202
rect 16452 7143 17942 7202
rect 18280 7143 19770 7202
rect 20108 7143 21598 7202
rect 0 6964 1490 7023
rect 1828 6964 3318 7023
rect 3656 6964 5146 7023
rect 5484 6964 6974 7023
rect 7312 6964 8802 7023
rect 9140 6964 10630 7023
rect 10968 6964 12458 7023
rect 12796 6964 14286 7023
rect 14624 6964 16114 7023
rect 16452 6964 17942 7023
rect 18280 6964 19770 7023
rect 20108 6964 21598 7023
rect 98 6952 128 6964
rect 290 6952 320 6964
rect 482 6952 512 6964
rect 674 6952 704 6964
rect 866 6952 896 6964
rect 1058 6952 1088 6964
rect 1250 6952 1280 6964
rect 1442 6952 1472 6964
rect 1926 6952 1956 6964
rect 2118 6952 2148 6964
rect 2310 6952 2340 6964
rect 2502 6952 2532 6964
rect 2694 6952 2724 6964
rect 2886 6952 2916 6964
rect 3078 6952 3108 6964
rect 3270 6952 3300 6964
rect 3754 6952 3784 6964
rect 3946 6952 3976 6964
rect 4138 6952 4168 6964
rect 4330 6952 4360 6964
rect 4522 6952 4552 6964
rect 4714 6952 4744 6964
rect 4906 6952 4936 6964
rect 5098 6952 5128 6964
rect 5582 6952 5612 6964
rect 5774 6952 5804 6964
rect 5966 6952 5996 6964
rect 6158 6952 6188 6964
rect 6350 6952 6380 6964
rect 6542 6952 6572 6964
rect 6734 6952 6764 6964
rect 6926 6952 6956 6964
rect 7410 6952 7440 6964
rect 7602 6952 7632 6964
rect 7794 6952 7824 6964
rect 7986 6952 8016 6964
rect 8178 6952 8208 6964
rect 8370 6952 8400 6964
rect 8562 6952 8592 6964
rect 8754 6952 8784 6964
rect 9238 6952 9268 6964
rect 9430 6952 9460 6964
rect 9622 6952 9652 6964
rect 9814 6952 9844 6964
rect 10006 6952 10036 6964
rect 10198 6952 10228 6964
rect 10390 6952 10420 6964
rect 10582 6952 10612 6964
rect 11066 6952 11096 6964
rect 11258 6952 11288 6964
rect 11450 6952 11480 6964
rect 11642 6952 11672 6964
rect 11834 6952 11864 6964
rect 12026 6952 12056 6964
rect 12218 6952 12248 6964
rect 12410 6952 12440 6964
rect 12894 6952 12924 6964
rect 13086 6952 13116 6964
rect 13278 6952 13308 6964
rect 13470 6952 13500 6964
rect 13662 6952 13692 6964
rect 13854 6952 13884 6964
rect 14046 6952 14076 6964
rect 14238 6952 14268 6964
rect 14722 6952 14752 6964
rect 14914 6952 14944 6964
rect 15106 6952 15136 6964
rect 15298 6952 15328 6964
rect 15490 6952 15520 6964
rect 15682 6952 15712 6964
rect 15874 6952 15904 6964
rect 16066 6952 16096 6964
rect 16550 6952 16580 6964
rect 16742 6952 16772 6964
rect 16934 6952 16964 6964
rect 17126 6952 17156 6964
rect 17318 6952 17348 6964
rect 17510 6952 17540 6964
rect 17702 6952 17732 6964
rect 17894 6952 17924 6964
rect 18378 6952 18408 6964
rect 18570 6952 18600 6964
rect 18762 6952 18792 6964
rect 18954 6952 18984 6964
rect 19146 6952 19176 6964
rect 19338 6952 19368 6964
rect 19530 6952 19560 6964
rect 19722 6952 19752 6964
rect 20206 6952 20236 6964
rect 20398 6952 20428 6964
rect 20590 6952 20620 6964
rect 20782 6952 20812 6964
rect 20974 6952 21004 6964
rect 21166 6952 21196 6964
rect 21358 6952 21388 6964
rect 21550 6952 21580 6964
rect 194 6488 224 6500
rect 386 6488 416 6500
rect 578 6488 608 6500
rect 770 6488 800 6500
rect 962 6488 992 6500
rect 1154 6488 1184 6500
rect 1346 6488 1376 6500
rect 2022 6488 2052 6500
rect 2214 6488 2244 6500
rect 2406 6488 2436 6500
rect 2598 6488 2628 6500
rect 2790 6488 2820 6500
rect 2982 6488 3012 6500
rect 3174 6488 3204 6500
rect 3850 6488 3880 6500
rect 4042 6488 4072 6500
rect 4234 6488 4264 6500
rect 4426 6488 4456 6500
rect 4618 6488 4648 6500
rect 4810 6488 4840 6500
rect 5002 6488 5032 6500
rect 5678 6488 5708 6500
rect 5870 6488 5900 6500
rect 6062 6488 6092 6500
rect 6254 6488 6284 6500
rect 6446 6488 6476 6500
rect 6638 6488 6668 6500
rect 6830 6488 6860 6500
rect 7506 6488 7536 6500
rect 7698 6488 7728 6500
rect 7890 6488 7920 6500
rect 8082 6488 8112 6500
rect 8274 6488 8304 6500
rect 8466 6488 8496 6500
rect 8658 6488 8688 6500
rect 9334 6488 9364 6500
rect 9526 6488 9556 6500
rect 9718 6488 9748 6500
rect 9910 6488 9940 6500
rect 10102 6488 10132 6500
rect 10294 6488 10324 6500
rect 10486 6488 10516 6500
rect 11162 6488 11192 6500
rect 11354 6488 11384 6500
rect 11546 6488 11576 6500
rect 11738 6488 11768 6500
rect 11930 6488 11960 6500
rect 12122 6488 12152 6500
rect 12314 6488 12344 6500
rect 12990 6488 13020 6500
rect 13182 6488 13212 6500
rect 13374 6488 13404 6500
rect 13566 6488 13596 6500
rect 13758 6488 13788 6500
rect 13950 6488 13980 6500
rect 14142 6488 14172 6500
rect 14818 6488 14848 6500
rect 15010 6488 15040 6500
rect 15202 6488 15232 6500
rect 15394 6488 15424 6500
rect 15586 6488 15616 6500
rect 15778 6488 15808 6500
rect 15970 6488 16000 6500
rect 16646 6488 16676 6500
rect 16838 6488 16868 6500
rect 17030 6488 17060 6500
rect 17222 6488 17252 6500
rect 17414 6488 17444 6500
rect 17606 6488 17636 6500
rect 17798 6488 17828 6500
rect 18474 6488 18504 6500
rect 18666 6488 18696 6500
rect 18858 6488 18888 6500
rect 19050 6488 19080 6500
rect 19242 6488 19272 6500
rect 19434 6488 19464 6500
rect 19626 6488 19656 6500
rect 20302 6488 20332 6500
rect 20494 6488 20524 6500
rect 20686 6488 20716 6500
rect 20878 6488 20908 6500
rect 21070 6488 21100 6500
rect 21262 6488 21292 6500
rect 21454 6488 21484 6500
rect 0 6429 1490 6488
rect 1828 6429 3318 6488
rect 3656 6429 5146 6488
rect 5484 6429 6974 6488
rect 7312 6429 8802 6488
rect 9140 6429 10630 6488
rect 10968 6429 12458 6488
rect 12796 6429 14286 6488
rect 14624 6429 16114 6488
rect 16452 6429 17942 6488
rect 18280 6429 19770 6488
rect 20108 6429 21598 6488
rect 0 6250 1490 6309
rect 1828 6250 3318 6309
rect 3656 6250 5146 6309
rect 5484 6250 6974 6309
rect 7312 6250 8802 6309
rect 9140 6250 10630 6309
rect 10968 6250 12458 6309
rect 12796 6250 14286 6309
rect 14624 6250 16114 6309
rect 16452 6250 17942 6309
rect 18280 6250 19770 6309
rect 20108 6250 21598 6309
rect 98 6238 128 6250
rect 290 6238 320 6250
rect 482 6238 512 6250
rect 674 6238 704 6250
rect 866 6238 896 6250
rect 1058 6238 1088 6250
rect 1250 6238 1280 6250
rect 1442 6238 1472 6250
rect 1926 6238 1956 6250
rect 2118 6238 2148 6250
rect 2310 6238 2340 6250
rect 2502 6238 2532 6250
rect 2694 6238 2724 6250
rect 2886 6238 2916 6250
rect 3078 6238 3108 6250
rect 3270 6238 3300 6250
rect 3754 6238 3784 6250
rect 3946 6238 3976 6250
rect 4138 6238 4168 6250
rect 4330 6238 4360 6250
rect 4522 6238 4552 6250
rect 4714 6238 4744 6250
rect 4906 6238 4936 6250
rect 5098 6238 5128 6250
rect 5582 6238 5612 6250
rect 5774 6238 5804 6250
rect 5966 6238 5996 6250
rect 6158 6238 6188 6250
rect 6350 6238 6380 6250
rect 6542 6238 6572 6250
rect 6734 6238 6764 6250
rect 6926 6238 6956 6250
rect 7410 6238 7440 6250
rect 7602 6238 7632 6250
rect 7794 6238 7824 6250
rect 7986 6238 8016 6250
rect 8178 6238 8208 6250
rect 8370 6238 8400 6250
rect 8562 6238 8592 6250
rect 8754 6238 8784 6250
rect 9238 6238 9268 6250
rect 9430 6238 9460 6250
rect 9622 6238 9652 6250
rect 9814 6238 9844 6250
rect 10006 6238 10036 6250
rect 10198 6238 10228 6250
rect 10390 6238 10420 6250
rect 10582 6238 10612 6250
rect 11066 6238 11096 6250
rect 11258 6238 11288 6250
rect 11450 6238 11480 6250
rect 11642 6238 11672 6250
rect 11834 6238 11864 6250
rect 12026 6238 12056 6250
rect 12218 6238 12248 6250
rect 12410 6238 12440 6250
rect 12894 6238 12924 6250
rect 13086 6238 13116 6250
rect 13278 6238 13308 6250
rect 13470 6238 13500 6250
rect 13662 6238 13692 6250
rect 13854 6238 13884 6250
rect 14046 6238 14076 6250
rect 14238 6238 14268 6250
rect 14722 6238 14752 6250
rect 14914 6238 14944 6250
rect 15106 6238 15136 6250
rect 15298 6238 15328 6250
rect 15490 6238 15520 6250
rect 15682 6238 15712 6250
rect 15874 6238 15904 6250
rect 16066 6238 16096 6250
rect 16550 6238 16580 6250
rect 16742 6238 16772 6250
rect 16934 6238 16964 6250
rect 17126 6238 17156 6250
rect 17318 6238 17348 6250
rect 17510 6238 17540 6250
rect 17702 6238 17732 6250
rect 17894 6238 17924 6250
rect 18378 6238 18408 6250
rect 18570 6238 18600 6250
rect 18762 6238 18792 6250
rect 18954 6238 18984 6250
rect 19146 6238 19176 6250
rect 19338 6238 19368 6250
rect 19530 6238 19560 6250
rect 19722 6238 19752 6250
rect 20206 6238 20236 6250
rect 20398 6238 20428 6250
rect 20590 6238 20620 6250
rect 20782 6238 20812 6250
rect 20974 6238 21004 6250
rect 21166 6238 21196 6250
rect 21358 6238 21388 6250
rect 21550 6238 21580 6250
rect 194 5774 224 5786
rect 386 5774 416 5786
rect 578 5774 608 5786
rect 770 5774 800 5786
rect 962 5774 992 5786
rect 1154 5774 1184 5786
rect 1346 5774 1376 5786
rect 2022 5774 2052 5786
rect 2214 5774 2244 5786
rect 2406 5774 2436 5786
rect 2598 5774 2628 5786
rect 2790 5774 2820 5786
rect 2982 5774 3012 5786
rect 3174 5774 3204 5786
rect 3850 5774 3880 5786
rect 4042 5774 4072 5786
rect 4234 5774 4264 5786
rect 4426 5774 4456 5786
rect 4618 5774 4648 5786
rect 4810 5774 4840 5786
rect 5002 5774 5032 5786
rect 5678 5774 5708 5786
rect 5870 5774 5900 5786
rect 6062 5774 6092 5786
rect 6254 5774 6284 5786
rect 6446 5774 6476 5786
rect 6638 5774 6668 5786
rect 6830 5774 6860 5786
rect 7506 5774 7536 5786
rect 7698 5774 7728 5786
rect 7890 5774 7920 5786
rect 8082 5774 8112 5786
rect 8274 5774 8304 5786
rect 8466 5774 8496 5786
rect 8658 5774 8688 5786
rect 9334 5774 9364 5786
rect 9526 5774 9556 5786
rect 9718 5774 9748 5786
rect 9910 5774 9940 5786
rect 10102 5774 10132 5786
rect 10294 5774 10324 5786
rect 10486 5774 10516 5786
rect 11162 5774 11192 5786
rect 11354 5774 11384 5786
rect 11546 5774 11576 5786
rect 11738 5774 11768 5786
rect 11930 5774 11960 5786
rect 12122 5774 12152 5786
rect 12314 5774 12344 5786
rect 12990 5774 13020 5786
rect 13182 5774 13212 5786
rect 13374 5774 13404 5786
rect 13566 5774 13596 5786
rect 13758 5774 13788 5786
rect 13950 5774 13980 5786
rect 14142 5774 14172 5786
rect 14818 5774 14848 5786
rect 15010 5774 15040 5786
rect 15202 5774 15232 5786
rect 15394 5774 15424 5786
rect 15586 5774 15616 5786
rect 15778 5774 15808 5786
rect 15970 5774 16000 5786
rect 16646 5774 16676 5786
rect 16838 5774 16868 5786
rect 17030 5774 17060 5786
rect 17222 5774 17252 5786
rect 17414 5774 17444 5786
rect 17606 5774 17636 5786
rect 17798 5774 17828 5786
rect 18474 5774 18504 5786
rect 18666 5774 18696 5786
rect 18858 5774 18888 5786
rect 19050 5774 19080 5786
rect 19242 5774 19272 5786
rect 19434 5774 19464 5786
rect 19626 5774 19656 5786
rect 20302 5774 20332 5786
rect 20494 5774 20524 5786
rect 20686 5774 20716 5786
rect 20878 5774 20908 5786
rect 21070 5774 21100 5786
rect 21262 5774 21292 5786
rect 21454 5774 21484 5786
rect 0 5715 1490 5774
rect 1828 5715 3318 5774
rect 3656 5715 5146 5774
rect 5484 5715 6974 5774
rect 7312 5715 8802 5774
rect 9140 5715 10630 5774
rect 10968 5715 12458 5774
rect 12796 5715 14286 5774
rect 14624 5715 16114 5774
rect 16452 5715 17942 5774
rect 18280 5715 19770 5774
rect 20108 5715 21598 5774
rect 0 5536 1490 5595
rect 1828 5536 3318 5595
rect 3656 5536 5146 5595
rect 5484 5536 6974 5595
rect 7312 5536 8802 5595
rect 9140 5536 10630 5595
rect 10968 5536 12458 5595
rect 12796 5536 14286 5595
rect 14624 5536 16114 5595
rect 16452 5536 17942 5595
rect 18280 5536 19770 5595
rect 20108 5536 21598 5595
rect 98 5524 128 5536
rect 290 5524 320 5536
rect 482 5524 512 5536
rect 674 5524 704 5536
rect 866 5524 896 5536
rect 1058 5524 1088 5536
rect 1250 5524 1280 5536
rect 1442 5524 1472 5536
rect 1926 5524 1956 5536
rect 2118 5524 2148 5536
rect 2310 5524 2340 5536
rect 2502 5524 2532 5536
rect 2694 5524 2724 5536
rect 2886 5524 2916 5536
rect 3078 5524 3108 5536
rect 3270 5524 3300 5536
rect 3754 5524 3784 5536
rect 3946 5524 3976 5536
rect 4138 5524 4168 5536
rect 4330 5524 4360 5536
rect 4522 5524 4552 5536
rect 4714 5524 4744 5536
rect 4906 5524 4936 5536
rect 5098 5524 5128 5536
rect 5582 5524 5612 5536
rect 5774 5524 5804 5536
rect 5966 5524 5996 5536
rect 6158 5524 6188 5536
rect 6350 5524 6380 5536
rect 6542 5524 6572 5536
rect 6734 5524 6764 5536
rect 6926 5524 6956 5536
rect 7410 5524 7440 5536
rect 7602 5524 7632 5536
rect 7794 5524 7824 5536
rect 7986 5524 8016 5536
rect 8178 5524 8208 5536
rect 8370 5524 8400 5536
rect 8562 5524 8592 5536
rect 8754 5524 8784 5536
rect 9238 5524 9268 5536
rect 9430 5524 9460 5536
rect 9622 5524 9652 5536
rect 9814 5524 9844 5536
rect 10006 5524 10036 5536
rect 10198 5524 10228 5536
rect 10390 5524 10420 5536
rect 10582 5524 10612 5536
rect 11066 5524 11096 5536
rect 11258 5524 11288 5536
rect 11450 5524 11480 5536
rect 11642 5524 11672 5536
rect 11834 5524 11864 5536
rect 12026 5524 12056 5536
rect 12218 5524 12248 5536
rect 12410 5524 12440 5536
rect 12894 5524 12924 5536
rect 13086 5524 13116 5536
rect 13278 5524 13308 5536
rect 13470 5524 13500 5536
rect 13662 5524 13692 5536
rect 13854 5524 13884 5536
rect 14046 5524 14076 5536
rect 14238 5524 14268 5536
rect 14722 5524 14752 5536
rect 14914 5524 14944 5536
rect 15106 5524 15136 5536
rect 15298 5524 15328 5536
rect 15490 5524 15520 5536
rect 15682 5524 15712 5536
rect 15874 5524 15904 5536
rect 16066 5524 16096 5536
rect 16550 5524 16580 5536
rect 16742 5524 16772 5536
rect 16934 5524 16964 5536
rect 17126 5524 17156 5536
rect 17318 5524 17348 5536
rect 17510 5524 17540 5536
rect 17702 5524 17732 5536
rect 17894 5524 17924 5536
rect 18378 5524 18408 5536
rect 18570 5524 18600 5536
rect 18762 5524 18792 5536
rect 18954 5524 18984 5536
rect 19146 5524 19176 5536
rect 19338 5524 19368 5536
rect 19530 5524 19560 5536
rect 19722 5524 19752 5536
rect 20206 5524 20236 5536
rect 20398 5524 20428 5536
rect 20590 5524 20620 5536
rect 20782 5524 20812 5536
rect 20974 5524 21004 5536
rect 21166 5524 21196 5536
rect 21358 5524 21388 5536
rect 21550 5524 21580 5536
rect 194 5060 224 5072
rect 386 5060 416 5072
rect 578 5060 608 5072
rect 770 5060 800 5072
rect 962 5060 992 5072
rect 1154 5060 1184 5072
rect 1346 5060 1376 5072
rect 2022 5060 2052 5072
rect 2214 5060 2244 5072
rect 2406 5060 2436 5072
rect 2598 5060 2628 5072
rect 2790 5060 2820 5072
rect 2982 5060 3012 5072
rect 3174 5060 3204 5072
rect 3850 5060 3880 5072
rect 4042 5060 4072 5072
rect 4234 5060 4264 5072
rect 4426 5060 4456 5072
rect 4618 5060 4648 5072
rect 4810 5060 4840 5072
rect 5002 5060 5032 5072
rect 5678 5060 5708 5072
rect 5870 5060 5900 5072
rect 6062 5060 6092 5072
rect 6254 5060 6284 5072
rect 6446 5060 6476 5072
rect 6638 5060 6668 5072
rect 6830 5060 6860 5072
rect 7506 5060 7536 5072
rect 7698 5060 7728 5072
rect 7890 5060 7920 5072
rect 8082 5060 8112 5072
rect 8274 5060 8304 5072
rect 8466 5060 8496 5072
rect 8658 5060 8688 5072
rect 9334 5060 9364 5072
rect 9526 5060 9556 5072
rect 9718 5060 9748 5072
rect 9910 5060 9940 5072
rect 10102 5060 10132 5072
rect 10294 5060 10324 5072
rect 10486 5060 10516 5072
rect 11162 5060 11192 5072
rect 11354 5060 11384 5072
rect 11546 5060 11576 5072
rect 11738 5060 11768 5072
rect 11930 5060 11960 5072
rect 12122 5060 12152 5072
rect 12314 5060 12344 5072
rect 12990 5060 13020 5072
rect 13182 5060 13212 5072
rect 13374 5060 13404 5072
rect 13566 5060 13596 5072
rect 13758 5060 13788 5072
rect 13950 5060 13980 5072
rect 14142 5060 14172 5072
rect 14818 5060 14848 5072
rect 15010 5060 15040 5072
rect 15202 5060 15232 5072
rect 15394 5060 15424 5072
rect 15586 5060 15616 5072
rect 15778 5060 15808 5072
rect 15970 5060 16000 5072
rect 16646 5060 16676 5072
rect 16838 5060 16868 5072
rect 17030 5060 17060 5072
rect 17222 5060 17252 5072
rect 17414 5060 17444 5072
rect 17606 5060 17636 5072
rect 17798 5060 17828 5072
rect 18474 5060 18504 5072
rect 18666 5060 18696 5072
rect 18858 5060 18888 5072
rect 19050 5060 19080 5072
rect 19242 5060 19272 5072
rect 19434 5060 19464 5072
rect 19626 5060 19656 5072
rect 20302 5060 20332 5072
rect 20494 5060 20524 5072
rect 20686 5060 20716 5072
rect 20878 5060 20908 5072
rect 21070 5060 21100 5072
rect 21262 5060 21292 5072
rect 21454 5060 21484 5072
rect 0 5001 1490 5060
rect 1828 5001 3318 5060
rect 3656 5001 5146 5060
rect 5484 5001 6974 5060
rect 7312 5001 8802 5060
rect 9140 5001 10630 5060
rect 10968 5001 12458 5060
rect 12796 5001 14286 5060
rect 14624 5001 16114 5060
rect 16452 5001 17942 5060
rect 18280 5001 19770 5060
rect 20108 5001 21598 5060
rect 0 4822 1490 4881
rect 1828 4822 3318 4881
rect 3656 4822 5146 4881
rect 5484 4822 6974 4881
rect 7312 4822 8802 4881
rect 9140 4822 10630 4881
rect 10968 4822 12458 4881
rect 12796 4822 14286 4881
rect 14624 4822 16114 4881
rect 16452 4822 17942 4881
rect 18280 4822 19770 4881
rect 20108 4822 21598 4881
rect 98 4810 128 4822
rect 290 4810 320 4822
rect 482 4810 512 4822
rect 674 4810 704 4822
rect 866 4810 896 4822
rect 1058 4810 1088 4822
rect 1250 4810 1280 4822
rect 1442 4810 1472 4822
rect 1926 4810 1956 4822
rect 2118 4810 2148 4822
rect 2310 4810 2340 4822
rect 2502 4810 2532 4822
rect 2694 4810 2724 4822
rect 2886 4810 2916 4822
rect 3078 4810 3108 4822
rect 3270 4810 3300 4822
rect 3754 4810 3784 4822
rect 3946 4810 3976 4822
rect 4138 4810 4168 4822
rect 4330 4810 4360 4822
rect 4522 4810 4552 4822
rect 4714 4810 4744 4822
rect 4906 4810 4936 4822
rect 5098 4810 5128 4822
rect 5582 4810 5612 4822
rect 5774 4810 5804 4822
rect 5966 4810 5996 4822
rect 6158 4810 6188 4822
rect 6350 4810 6380 4822
rect 6542 4810 6572 4822
rect 6734 4810 6764 4822
rect 6926 4810 6956 4822
rect 7410 4810 7440 4822
rect 7602 4810 7632 4822
rect 7794 4810 7824 4822
rect 7986 4810 8016 4822
rect 8178 4810 8208 4822
rect 8370 4810 8400 4822
rect 8562 4810 8592 4822
rect 8754 4810 8784 4822
rect 9238 4810 9268 4822
rect 9430 4810 9460 4822
rect 9622 4810 9652 4822
rect 9814 4810 9844 4822
rect 10006 4810 10036 4822
rect 10198 4810 10228 4822
rect 10390 4810 10420 4822
rect 10582 4810 10612 4822
rect 11066 4810 11096 4822
rect 11258 4810 11288 4822
rect 11450 4810 11480 4822
rect 11642 4810 11672 4822
rect 11834 4810 11864 4822
rect 12026 4810 12056 4822
rect 12218 4810 12248 4822
rect 12410 4810 12440 4822
rect 12894 4810 12924 4822
rect 13086 4810 13116 4822
rect 13278 4810 13308 4822
rect 13470 4810 13500 4822
rect 13662 4810 13692 4822
rect 13854 4810 13884 4822
rect 14046 4810 14076 4822
rect 14238 4810 14268 4822
rect 14722 4810 14752 4822
rect 14914 4810 14944 4822
rect 15106 4810 15136 4822
rect 15298 4810 15328 4822
rect 15490 4810 15520 4822
rect 15682 4810 15712 4822
rect 15874 4810 15904 4822
rect 16066 4810 16096 4822
rect 16550 4810 16580 4822
rect 16742 4810 16772 4822
rect 16934 4810 16964 4822
rect 17126 4810 17156 4822
rect 17318 4810 17348 4822
rect 17510 4810 17540 4822
rect 17702 4810 17732 4822
rect 17894 4810 17924 4822
rect 18378 4810 18408 4822
rect 18570 4810 18600 4822
rect 18762 4810 18792 4822
rect 18954 4810 18984 4822
rect 19146 4810 19176 4822
rect 19338 4810 19368 4822
rect 19530 4810 19560 4822
rect 19722 4810 19752 4822
rect 20206 4810 20236 4822
rect 20398 4810 20428 4822
rect 20590 4810 20620 4822
rect 20782 4810 20812 4822
rect 20974 4810 21004 4822
rect 21166 4810 21196 4822
rect 21358 4810 21388 4822
rect 21550 4810 21580 4822
rect 194 4346 224 4358
rect 386 4346 416 4358
rect 578 4346 608 4358
rect 770 4346 800 4358
rect 962 4346 992 4358
rect 1154 4346 1184 4358
rect 1346 4346 1376 4358
rect 2022 4346 2052 4358
rect 2214 4346 2244 4358
rect 2406 4346 2436 4358
rect 2598 4346 2628 4358
rect 2790 4346 2820 4358
rect 2982 4346 3012 4358
rect 3174 4346 3204 4358
rect 3850 4346 3880 4358
rect 4042 4346 4072 4358
rect 4234 4346 4264 4358
rect 4426 4346 4456 4358
rect 4618 4346 4648 4358
rect 4810 4346 4840 4358
rect 5002 4346 5032 4358
rect 5678 4346 5708 4358
rect 5870 4346 5900 4358
rect 6062 4346 6092 4358
rect 6254 4346 6284 4358
rect 6446 4346 6476 4358
rect 6638 4346 6668 4358
rect 6830 4346 6860 4358
rect 7506 4346 7536 4358
rect 7698 4346 7728 4358
rect 7890 4346 7920 4358
rect 8082 4346 8112 4358
rect 8274 4346 8304 4358
rect 8466 4346 8496 4358
rect 8658 4346 8688 4358
rect 9334 4346 9364 4358
rect 9526 4346 9556 4358
rect 9718 4346 9748 4358
rect 9910 4346 9940 4358
rect 10102 4346 10132 4358
rect 10294 4346 10324 4358
rect 10486 4346 10516 4358
rect 11162 4346 11192 4358
rect 11354 4346 11384 4358
rect 11546 4346 11576 4358
rect 11738 4346 11768 4358
rect 11930 4346 11960 4358
rect 12122 4346 12152 4358
rect 12314 4346 12344 4358
rect 12990 4346 13020 4358
rect 13182 4346 13212 4358
rect 13374 4346 13404 4358
rect 13566 4346 13596 4358
rect 13758 4346 13788 4358
rect 13950 4346 13980 4358
rect 14142 4346 14172 4358
rect 14818 4346 14848 4358
rect 15010 4346 15040 4358
rect 15202 4346 15232 4358
rect 15394 4346 15424 4358
rect 15586 4346 15616 4358
rect 15778 4346 15808 4358
rect 15970 4346 16000 4358
rect 16646 4346 16676 4358
rect 16838 4346 16868 4358
rect 17030 4346 17060 4358
rect 17222 4346 17252 4358
rect 17414 4346 17444 4358
rect 17606 4346 17636 4358
rect 17798 4346 17828 4358
rect 18474 4346 18504 4358
rect 18666 4346 18696 4358
rect 18858 4346 18888 4358
rect 19050 4346 19080 4358
rect 19242 4346 19272 4358
rect 19434 4346 19464 4358
rect 19626 4346 19656 4358
rect 20302 4346 20332 4358
rect 20494 4346 20524 4358
rect 20686 4346 20716 4358
rect 20878 4346 20908 4358
rect 21070 4346 21100 4358
rect 21262 4346 21292 4358
rect 21454 4346 21484 4358
rect 0 4287 1490 4346
rect 1828 4287 3318 4346
rect 3656 4287 5146 4346
rect 5484 4287 6974 4346
rect 7312 4287 8802 4346
rect 9140 4287 10630 4346
rect 10968 4287 12458 4346
rect 12796 4287 14286 4346
rect 14624 4287 16114 4346
rect 16452 4287 17942 4346
rect 18280 4287 19770 4346
rect 20108 4287 21598 4346
rect 0 4108 1490 4167
rect 1828 4108 3318 4167
rect 3656 4108 5146 4167
rect 5484 4108 6974 4167
rect 7312 4108 8802 4167
rect 9140 4108 10630 4167
rect 10968 4108 12458 4167
rect 12796 4108 14286 4167
rect 14624 4108 16114 4167
rect 16452 4108 17942 4167
rect 18280 4108 19770 4167
rect 20108 4108 21598 4167
rect 98 4096 128 4108
rect 290 4096 320 4108
rect 482 4096 512 4108
rect 674 4096 704 4108
rect 866 4096 896 4108
rect 1058 4096 1088 4108
rect 1250 4096 1280 4108
rect 1442 4096 1472 4108
rect 1926 4096 1956 4108
rect 2118 4096 2148 4108
rect 2310 4096 2340 4108
rect 2502 4096 2532 4108
rect 2694 4096 2724 4108
rect 2886 4096 2916 4108
rect 3078 4096 3108 4108
rect 3270 4096 3300 4108
rect 3754 4096 3784 4108
rect 3946 4096 3976 4108
rect 4138 4096 4168 4108
rect 4330 4096 4360 4108
rect 4522 4096 4552 4108
rect 4714 4096 4744 4108
rect 4906 4096 4936 4108
rect 5098 4096 5128 4108
rect 5582 4096 5612 4108
rect 5774 4096 5804 4108
rect 5966 4096 5996 4108
rect 6158 4096 6188 4108
rect 6350 4096 6380 4108
rect 6542 4096 6572 4108
rect 6734 4096 6764 4108
rect 6926 4096 6956 4108
rect 7410 4096 7440 4108
rect 7602 4096 7632 4108
rect 7794 4096 7824 4108
rect 7986 4096 8016 4108
rect 8178 4096 8208 4108
rect 8370 4096 8400 4108
rect 8562 4096 8592 4108
rect 8754 4096 8784 4108
rect 9238 4096 9268 4108
rect 9430 4096 9460 4108
rect 9622 4096 9652 4108
rect 9814 4096 9844 4108
rect 10006 4096 10036 4108
rect 10198 4096 10228 4108
rect 10390 4096 10420 4108
rect 10582 4096 10612 4108
rect 11066 4096 11096 4108
rect 11258 4096 11288 4108
rect 11450 4096 11480 4108
rect 11642 4096 11672 4108
rect 11834 4096 11864 4108
rect 12026 4096 12056 4108
rect 12218 4096 12248 4108
rect 12410 4096 12440 4108
rect 12894 4096 12924 4108
rect 13086 4096 13116 4108
rect 13278 4096 13308 4108
rect 13470 4096 13500 4108
rect 13662 4096 13692 4108
rect 13854 4096 13884 4108
rect 14046 4096 14076 4108
rect 14238 4096 14268 4108
rect 14722 4096 14752 4108
rect 14914 4096 14944 4108
rect 15106 4096 15136 4108
rect 15298 4096 15328 4108
rect 15490 4096 15520 4108
rect 15682 4096 15712 4108
rect 15874 4096 15904 4108
rect 16066 4096 16096 4108
rect 16550 4096 16580 4108
rect 16742 4096 16772 4108
rect 16934 4096 16964 4108
rect 17126 4096 17156 4108
rect 17318 4096 17348 4108
rect 17510 4096 17540 4108
rect 17702 4096 17732 4108
rect 17894 4096 17924 4108
rect 18378 4096 18408 4108
rect 18570 4096 18600 4108
rect 18762 4096 18792 4108
rect 18954 4096 18984 4108
rect 19146 4096 19176 4108
rect 19338 4096 19368 4108
rect 19530 4096 19560 4108
rect 19722 4096 19752 4108
rect 20206 4096 20236 4108
rect 20398 4096 20428 4108
rect 20590 4096 20620 4108
rect 20782 4096 20812 4108
rect 20974 4096 21004 4108
rect 21166 4096 21196 4108
rect 21358 4096 21388 4108
rect 21550 4096 21580 4108
rect 194 3632 224 3644
rect 386 3632 416 3644
rect 578 3632 608 3644
rect 770 3632 800 3644
rect 962 3632 992 3644
rect 1154 3632 1184 3644
rect 1346 3632 1376 3644
rect 2022 3632 2052 3644
rect 2214 3632 2244 3644
rect 2406 3632 2436 3644
rect 2598 3632 2628 3644
rect 2790 3632 2820 3644
rect 2982 3632 3012 3644
rect 3174 3632 3204 3644
rect 3850 3632 3880 3644
rect 4042 3632 4072 3644
rect 4234 3632 4264 3644
rect 4426 3632 4456 3644
rect 4618 3632 4648 3644
rect 4810 3632 4840 3644
rect 5002 3632 5032 3644
rect 5678 3632 5708 3644
rect 5870 3632 5900 3644
rect 6062 3632 6092 3644
rect 6254 3632 6284 3644
rect 6446 3632 6476 3644
rect 6638 3632 6668 3644
rect 6830 3632 6860 3644
rect 7506 3632 7536 3644
rect 7698 3632 7728 3644
rect 7890 3632 7920 3644
rect 8082 3632 8112 3644
rect 8274 3632 8304 3644
rect 8466 3632 8496 3644
rect 8658 3632 8688 3644
rect 9334 3632 9364 3644
rect 9526 3632 9556 3644
rect 9718 3632 9748 3644
rect 9910 3632 9940 3644
rect 10102 3632 10132 3644
rect 10294 3632 10324 3644
rect 10486 3632 10516 3644
rect 11162 3632 11192 3644
rect 11354 3632 11384 3644
rect 11546 3632 11576 3644
rect 11738 3632 11768 3644
rect 11930 3632 11960 3644
rect 12122 3632 12152 3644
rect 12314 3632 12344 3644
rect 12990 3632 13020 3644
rect 13182 3632 13212 3644
rect 13374 3632 13404 3644
rect 13566 3632 13596 3644
rect 13758 3632 13788 3644
rect 13950 3632 13980 3644
rect 14142 3632 14172 3644
rect 14818 3632 14848 3644
rect 15010 3632 15040 3644
rect 15202 3632 15232 3644
rect 15394 3632 15424 3644
rect 15586 3632 15616 3644
rect 15778 3632 15808 3644
rect 15970 3632 16000 3644
rect 16646 3632 16676 3644
rect 16838 3632 16868 3644
rect 17030 3632 17060 3644
rect 17222 3632 17252 3644
rect 17414 3632 17444 3644
rect 17606 3632 17636 3644
rect 17798 3632 17828 3644
rect 18474 3632 18504 3644
rect 18666 3632 18696 3644
rect 18858 3632 18888 3644
rect 19050 3632 19080 3644
rect 19242 3632 19272 3644
rect 19434 3632 19464 3644
rect 19626 3632 19656 3644
rect 20302 3632 20332 3644
rect 20494 3632 20524 3644
rect 20686 3632 20716 3644
rect 20878 3632 20908 3644
rect 21070 3632 21100 3644
rect 21262 3632 21292 3644
rect 21454 3632 21484 3644
rect 0 3573 1490 3632
rect 1828 3573 3318 3632
rect 3656 3573 5146 3632
rect 5484 3573 6974 3632
rect 7312 3573 8802 3632
rect 9140 3573 10630 3632
rect 10968 3573 12458 3632
rect 12796 3573 14286 3632
rect 14624 3573 16114 3632
rect 16452 3573 17942 3632
rect 18280 3573 19770 3632
rect 20108 3573 21598 3632
rect 0 3394 1490 3453
rect 1828 3394 3318 3453
rect 3656 3394 5146 3453
rect 5484 3394 6974 3453
rect 7312 3394 8802 3453
rect 9140 3394 10630 3453
rect 10968 3394 12458 3453
rect 12796 3394 14286 3453
rect 14624 3394 16114 3453
rect 16452 3394 17942 3453
rect 18280 3394 19770 3453
rect 20108 3394 21598 3453
rect 98 3382 128 3394
rect 290 3382 320 3394
rect 482 3382 512 3394
rect 674 3382 704 3394
rect 866 3382 896 3394
rect 1058 3382 1088 3394
rect 1250 3382 1280 3394
rect 1442 3382 1472 3394
rect 1926 3382 1956 3394
rect 2118 3382 2148 3394
rect 2310 3382 2340 3394
rect 2502 3382 2532 3394
rect 2694 3382 2724 3394
rect 2886 3382 2916 3394
rect 3078 3382 3108 3394
rect 3270 3382 3300 3394
rect 3754 3382 3784 3394
rect 3946 3382 3976 3394
rect 4138 3382 4168 3394
rect 4330 3382 4360 3394
rect 4522 3382 4552 3394
rect 4714 3382 4744 3394
rect 4906 3382 4936 3394
rect 5098 3382 5128 3394
rect 5582 3382 5612 3394
rect 5774 3382 5804 3394
rect 5966 3382 5996 3394
rect 6158 3382 6188 3394
rect 6350 3382 6380 3394
rect 6542 3382 6572 3394
rect 6734 3382 6764 3394
rect 6926 3382 6956 3394
rect 7410 3382 7440 3394
rect 7602 3382 7632 3394
rect 7794 3382 7824 3394
rect 7986 3382 8016 3394
rect 8178 3382 8208 3394
rect 8370 3382 8400 3394
rect 8562 3382 8592 3394
rect 8754 3382 8784 3394
rect 9238 3382 9268 3394
rect 9430 3382 9460 3394
rect 9622 3382 9652 3394
rect 9814 3382 9844 3394
rect 10006 3382 10036 3394
rect 10198 3382 10228 3394
rect 10390 3382 10420 3394
rect 10582 3382 10612 3394
rect 11066 3382 11096 3394
rect 11258 3382 11288 3394
rect 11450 3382 11480 3394
rect 11642 3382 11672 3394
rect 11834 3382 11864 3394
rect 12026 3382 12056 3394
rect 12218 3382 12248 3394
rect 12410 3382 12440 3394
rect 12894 3382 12924 3394
rect 13086 3382 13116 3394
rect 13278 3382 13308 3394
rect 13470 3382 13500 3394
rect 13662 3382 13692 3394
rect 13854 3382 13884 3394
rect 14046 3382 14076 3394
rect 14238 3382 14268 3394
rect 14722 3382 14752 3394
rect 14914 3382 14944 3394
rect 15106 3382 15136 3394
rect 15298 3382 15328 3394
rect 15490 3382 15520 3394
rect 15682 3382 15712 3394
rect 15874 3382 15904 3394
rect 16066 3382 16096 3394
rect 16550 3382 16580 3394
rect 16742 3382 16772 3394
rect 16934 3382 16964 3394
rect 17126 3382 17156 3394
rect 17318 3382 17348 3394
rect 17510 3382 17540 3394
rect 17702 3382 17732 3394
rect 17894 3382 17924 3394
rect 18378 3382 18408 3394
rect 18570 3382 18600 3394
rect 18762 3382 18792 3394
rect 18954 3382 18984 3394
rect 19146 3382 19176 3394
rect 19338 3382 19368 3394
rect 19530 3382 19560 3394
rect 19722 3382 19752 3394
rect 20206 3382 20236 3394
rect 20398 3382 20428 3394
rect 20590 3382 20620 3394
rect 20782 3382 20812 3394
rect 20974 3382 21004 3394
rect 21166 3382 21196 3394
rect 21358 3382 21388 3394
rect 21550 3382 21580 3394
rect 194 2918 224 2930
rect 386 2918 416 2930
rect 578 2918 608 2930
rect 770 2918 800 2930
rect 962 2918 992 2930
rect 1154 2918 1184 2930
rect 1346 2918 1376 2930
rect 2022 2918 2052 2930
rect 2214 2918 2244 2930
rect 2406 2918 2436 2930
rect 2598 2918 2628 2930
rect 2790 2918 2820 2930
rect 2982 2918 3012 2930
rect 3174 2918 3204 2930
rect 3850 2918 3880 2930
rect 4042 2918 4072 2930
rect 4234 2918 4264 2930
rect 4426 2918 4456 2930
rect 4618 2918 4648 2930
rect 4810 2918 4840 2930
rect 5002 2918 5032 2930
rect 5678 2918 5708 2930
rect 5870 2918 5900 2930
rect 6062 2918 6092 2930
rect 6254 2918 6284 2930
rect 6446 2918 6476 2930
rect 6638 2918 6668 2930
rect 6830 2918 6860 2930
rect 7506 2918 7536 2930
rect 7698 2918 7728 2930
rect 7890 2918 7920 2930
rect 8082 2918 8112 2930
rect 8274 2918 8304 2930
rect 8466 2918 8496 2930
rect 8658 2918 8688 2930
rect 9334 2918 9364 2930
rect 9526 2918 9556 2930
rect 9718 2918 9748 2930
rect 9910 2918 9940 2930
rect 10102 2918 10132 2930
rect 10294 2918 10324 2930
rect 10486 2918 10516 2930
rect 11162 2918 11192 2930
rect 11354 2918 11384 2930
rect 11546 2918 11576 2930
rect 11738 2918 11768 2930
rect 11930 2918 11960 2930
rect 12122 2918 12152 2930
rect 12314 2918 12344 2930
rect 12990 2918 13020 2930
rect 13182 2918 13212 2930
rect 13374 2918 13404 2930
rect 13566 2918 13596 2930
rect 13758 2918 13788 2930
rect 13950 2918 13980 2930
rect 14142 2918 14172 2930
rect 14818 2918 14848 2930
rect 15010 2918 15040 2930
rect 15202 2918 15232 2930
rect 15394 2918 15424 2930
rect 15586 2918 15616 2930
rect 15778 2918 15808 2930
rect 15970 2918 16000 2930
rect 16646 2918 16676 2930
rect 16838 2918 16868 2930
rect 17030 2918 17060 2930
rect 17222 2918 17252 2930
rect 17414 2918 17444 2930
rect 17606 2918 17636 2930
rect 17798 2918 17828 2930
rect 18474 2918 18504 2930
rect 18666 2918 18696 2930
rect 18858 2918 18888 2930
rect 19050 2918 19080 2930
rect 19242 2918 19272 2930
rect 19434 2918 19464 2930
rect 19626 2918 19656 2930
rect 20302 2918 20332 2930
rect 20494 2918 20524 2930
rect 20686 2918 20716 2930
rect 20878 2918 20908 2930
rect 21070 2918 21100 2930
rect 21262 2918 21292 2930
rect 21454 2918 21484 2930
rect 0 2859 1490 2918
rect 1828 2859 3318 2918
rect 3656 2859 5146 2918
rect 5484 2859 6974 2918
rect 7312 2859 8802 2918
rect 9140 2859 10630 2918
rect 10968 2859 12458 2918
rect 12796 2859 14286 2918
rect 14624 2859 16114 2918
rect 16452 2859 17942 2918
rect 18280 2859 19770 2918
rect 20108 2859 21598 2918
rect 0 2680 1490 2739
rect 1828 2680 3318 2739
rect 3656 2680 5146 2739
rect 5484 2680 6974 2739
rect 7312 2680 8802 2739
rect 9140 2680 10630 2739
rect 10968 2680 12458 2739
rect 12796 2680 14286 2739
rect 14624 2680 16114 2739
rect 16452 2680 17942 2739
rect 18280 2680 19770 2739
rect 20108 2680 21598 2739
rect 98 2668 128 2680
rect 290 2668 320 2680
rect 482 2668 512 2680
rect 674 2668 704 2680
rect 866 2668 896 2680
rect 1058 2668 1088 2680
rect 1250 2668 1280 2680
rect 1442 2668 1472 2680
rect 1926 2668 1956 2680
rect 2118 2668 2148 2680
rect 2310 2668 2340 2680
rect 2502 2668 2532 2680
rect 2694 2668 2724 2680
rect 2886 2668 2916 2680
rect 3078 2668 3108 2680
rect 3270 2668 3300 2680
rect 3754 2668 3784 2680
rect 3946 2668 3976 2680
rect 4138 2668 4168 2680
rect 4330 2668 4360 2680
rect 4522 2668 4552 2680
rect 4714 2668 4744 2680
rect 4906 2668 4936 2680
rect 5098 2668 5128 2680
rect 5582 2668 5612 2680
rect 5774 2668 5804 2680
rect 5966 2668 5996 2680
rect 6158 2668 6188 2680
rect 6350 2668 6380 2680
rect 6542 2668 6572 2680
rect 6734 2668 6764 2680
rect 6926 2668 6956 2680
rect 7410 2668 7440 2680
rect 7602 2668 7632 2680
rect 7794 2668 7824 2680
rect 7986 2668 8016 2680
rect 8178 2668 8208 2680
rect 8370 2668 8400 2680
rect 8562 2668 8592 2680
rect 8754 2668 8784 2680
rect 9238 2668 9268 2680
rect 9430 2668 9460 2680
rect 9622 2668 9652 2680
rect 9814 2668 9844 2680
rect 10006 2668 10036 2680
rect 10198 2668 10228 2680
rect 10390 2668 10420 2680
rect 10582 2668 10612 2680
rect 11066 2668 11096 2680
rect 11258 2668 11288 2680
rect 11450 2668 11480 2680
rect 11642 2668 11672 2680
rect 11834 2668 11864 2680
rect 12026 2668 12056 2680
rect 12218 2668 12248 2680
rect 12410 2668 12440 2680
rect 12894 2668 12924 2680
rect 13086 2668 13116 2680
rect 13278 2668 13308 2680
rect 13470 2668 13500 2680
rect 13662 2668 13692 2680
rect 13854 2668 13884 2680
rect 14046 2668 14076 2680
rect 14238 2668 14268 2680
rect 14722 2668 14752 2680
rect 14914 2668 14944 2680
rect 15106 2668 15136 2680
rect 15298 2668 15328 2680
rect 15490 2668 15520 2680
rect 15682 2668 15712 2680
rect 15874 2668 15904 2680
rect 16066 2668 16096 2680
rect 16550 2668 16580 2680
rect 16742 2668 16772 2680
rect 16934 2668 16964 2680
rect 17126 2668 17156 2680
rect 17318 2668 17348 2680
rect 17510 2668 17540 2680
rect 17702 2668 17732 2680
rect 17894 2668 17924 2680
rect 18378 2668 18408 2680
rect 18570 2668 18600 2680
rect 18762 2668 18792 2680
rect 18954 2668 18984 2680
rect 19146 2668 19176 2680
rect 19338 2668 19368 2680
rect 19530 2668 19560 2680
rect 19722 2668 19752 2680
rect 20206 2668 20236 2680
rect 20398 2668 20428 2680
rect 20590 2668 20620 2680
rect 20782 2668 20812 2680
rect 20974 2668 21004 2680
rect 21166 2668 21196 2680
rect 21358 2668 21388 2680
rect 21550 2668 21580 2680
rect 194 2204 224 2216
rect 386 2204 416 2216
rect 578 2204 608 2216
rect 770 2204 800 2216
rect 962 2204 992 2216
rect 1154 2204 1184 2216
rect 1346 2204 1376 2216
rect 2022 2204 2052 2216
rect 2214 2204 2244 2216
rect 2406 2204 2436 2216
rect 2598 2204 2628 2216
rect 2790 2204 2820 2216
rect 2982 2204 3012 2216
rect 3174 2204 3204 2216
rect 3850 2204 3880 2216
rect 4042 2204 4072 2216
rect 4234 2204 4264 2216
rect 4426 2204 4456 2216
rect 4618 2204 4648 2216
rect 4810 2204 4840 2216
rect 5002 2204 5032 2216
rect 5678 2204 5708 2216
rect 5870 2204 5900 2216
rect 6062 2204 6092 2216
rect 6254 2204 6284 2216
rect 6446 2204 6476 2216
rect 6638 2204 6668 2216
rect 6830 2204 6860 2216
rect 7506 2204 7536 2216
rect 7698 2204 7728 2216
rect 7890 2204 7920 2216
rect 8082 2204 8112 2216
rect 8274 2204 8304 2216
rect 8466 2204 8496 2216
rect 8658 2204 8688 2216
rect 9334 2204 9364 2216
rect 9526 2204 9556 2216
rect 9718 2204 9748 2216
rect 9910 2204 9940 2216
rect 10102 2204 10132 2216
rect 10294 2204 10324 2216
rect 10486 2204 10516 2216
rect 11162 2204 11192 2216
rect 11354 2204 11384 2216
rect 11546 2204 11576 2216
rect 11738 2204 11768 2216
rect 11930 2204 11960 2216
rect 12122 2204 12152 2216
rect 12314 2204 12344 2216
rect 12990 2204 13020 2216
rect 13182 2204 13212 2216
rect 13374 2204 13404 2216
rect 13566 2204 13596 2216
rect 13758 2204 13788 2216
rect 13950 2204 13980 2216
rect 14142 2204 14172 2216
rect 14818 2204 14848 2216
rect 15010 2204 15040 2216
rect 15202 2204 15232 2216
rect 15394 2204 15424 2216
rect 15586 2204 15616 2216
rect 15778 2204 15808 2216
rect 15970 2204 16000 2216
rect 16646 2204 16676 2216
rect 16838 2204 16868 2216
rect 17030 2204 17060 2216
rect 17222 2204 17252 2216
rect 17414 2204 17444 2216
rect 17606 2204 17636 2216
rect 17798 2204 17828 2216
rect 18474 2204 18504 2216
rect 18666 2204 18696 2216
rect 18858 2204 18888 2216
rect 19050 2204 19080 2216
rect 19242 2204 19272 2216
rect 19434 2204 19464 2216
rect 19626 2204 19656 2216
rect 20302 2204 20332 2216
rect 20494 2204 20524 2216
rect 20686 2204 20716 2216
rect 20878 2204 20908 2216
rect 21070 2204 21100 2216
rect 21262 2204 21292 2216
rect 21454 2204 21484 2216
rect 0 2145 1490 2204
rect 1828 2145 3318 2204
rect 3656 2145 5146 2204
rect 5484 2145 6974 2204
rect 7312 2145 8802 2204
rect 9140 2145 10630 2204
rect 10968 2145 12458 2204
rect 12796 2145 14286 2204
rect 14624 2145 16114 2204
rect 16452 2145 17942 2204
rect 18280 2145 19770 2204
rect 20108 2145 21598 2204
rect 0 1966 1490 2025
rect 1828 1966 3318 2025
rect 3656 1966 5146 2025
rect 5484 1966 6974 2025
rect 7312 1966 8802 2025
rect 9140 1966 10630 2025
rect 10968 1966 12458 2025
rect 12796 1966 14286 2025
rect 14624 1966 16114 2025
rect 16452 1966 17942 2025
rect 18280 1966 19770 2025
rect 20108 1966 21598 2025
rect 98 1954 128 1966
rect 290 1954 320 1966
rect 482 1954 512 1966
rect 674 1954 704 1966
rect 866 1954 896 1966
rect 1058 1954 1088 1966
rect 1250 1954 1280 1966
rect 1442 1954 1472 1966
rect 1926 1954 1956 1966
rect 2118 1954 2148 1966
rect 2310 1954 2340 1966
rect 2502 1954 2532 1966
rect 2694 1954 2724 1966
rect 2886 1954 2916 1966
rect 3078 1954 3108 1966
rect 3270 1954 3300 1966
rect 3754 1954 3784 1966
rect 3946 1954 3976 1966
rect 4138 1954 4168 1966
rect 4330 1954 4360 1966
rect 4522 1954 4552 1966
rect 4714 1954 4744 1966
rect 4906 1954 4936 1966
rect 5098 1954 5128 1966
rect 5582 1954 5612 1966
rect 5774 1954 5804 1966
rect 5966 1954 5996 1966
rect 6158 1954 6188 1966
rect 6350 1954 6380 1966
rect 6542 1954 6572 1966
rect 6734 1954 6764 1966
rect 6926 1954 6956 1966
rect 7410 1954 7440 1966
rect 7602 1954 7632 1966
rect 7794 1954 7824 1966
rect 7986 1954 8016 1966
rect 8178 1954 8208 1966
rect 8370 1954 8400 1966
rect 8562 1954 8592 1966
rect 8754 1954 8784 1966
rect 9238 1954 9268 1966
rect 9430 1954 9460 1966
rect 9622 1954 9652 1966
rect 9814 1954 9844 1966
rect 10006 1954 10036 1966
rect 10198 1954 10228 1966
rect 10390 1954 10420 1966
rect 10582 1954 10612 1966
rect 11066 1954 11096 1966
rect 11258 1954 11288 1966
rect 11450 1954 11480 1966
rect 11642 1954 11672 1966
rect 11834 1954 11864 1966
rect 12026 1954 12056 1966
rect 12218 1954 12248 1966
rect 12410 1954 12440 1966
rect 12894 1954 12924 1966
rect 13086 1954 13116 1966
rect 13278 1954 13308 1966
rect 13470 1954 13500 1966
rect 13662 1954 13692 1966
rect 13854 1954 13884 1966
rect 14046 1954 14076 1966
rect 14238 1954 14268 1966
rect 14722 1954 14752 1966
rect 14914 1954 14944 1966
rect 15106 1954 15136 1966
rect 15298 1954 15328 1966
rect 15490 1954 15520 1966
rect 15682 1954 15712 1966
rect 15874 1954 15904 1966
rect 16066 1954 16096 1966
rect 16550 1954 16580 1966
rect 16742 1954 16772 1966
rect 16934 1954 16964 1966
rect 17126 1954 17156 1966
rect 17318 1954 17348 1966
rect 17510 1954 17540 1966
rect 17702 1954 17732 1966
rect 17894 1954 17924 1966
rect 18378 1954 18408 1966
rect 18570 1954 18600 1966
rect 18762 1954 18792 1966
rect 18954 1954 18984 1966
rect 19146 1954 19176 1966
rect 19338 1954 19368 1966
rect 19530 1954 19560 1966
rect 19722 1954 19752 1966
rect 20206 1954 20236 1966
rect 20398 1954 20428 1966
rect 20590 1954 20620 1966
rect 20782 1954 20812 1966
rect 20974 1954 21004 1966
rect 21166 1954 21196 1966
rect 21358 1954 21388 1966
rect 21550 1954 21580 1966
rect 194 1490 224 1502
rect 386 1490 416 1502
rect 578 1490 608 1502
rect 770 1490 800 1502
rect 962 1490 992 1502
rect 1154 1490 1184 1502
rect 1346 1490 1376 1502
rect 2022 1490 2052 1502
rect 2214 1490 2244 1502
rect 2406 1490 2436 1502
rect 2598 1490 2628 1502
rect 2790 1490 2820 1502
rect 2982 1490 3012 1502
rect 3174 1490 3204 1502
rect 3850 1490 3880 1502
rect 4042 1490 4072 1502
rect 4234 1490 4264 1502
rect 4426 1490 4456 1502
rect 4618 1490 4648 1502
rect 4810 1490 4840 1502
rect 5002 1490 5032 1502
rect 5678 1490 5708 1502
rect 5870 1490 5900 1502
rect 6062 1490 6092 1502
rect 6254 1490 6284 1502
rect 6446 1490 6476 1502
rect 6638 1490 6668 1502
rect 6830 1490 6860 1502
rect 7506 1490 7536 1502
rect 7698 1490 7728 1502
rect 7890 1490 7920 1502
rect 8082 1490 8112 1502
rect 8274 1490 8304 1502
rect 8466 1490 8496 1502
rect 8658 1490 8688 1502
rect 9334 1490 9364 1502
rect 9526 1490 9556 1502
rect 9718 1490 9748 1502
rect 9910 1490 9940 1502
rect 10102 1490 10132 1502
rect 10294 1490 10324 1502
rect 10486 1490 10516 1502
rect 11162 1490 11192 1502
rect 11354 1490 11384 1502
rect 11546 1490 11576 1502
rect 11738 1490 11768 1502
rect 11930 1490 11960 1502
rect 12122 1490 12152 1502
rect 12314 1490 12344 1502
rect 12990 1490 13020 1502
rect 13182 1490 13212 1502
rect 13374 1490 13404 1502
rect 13566 1490 13596 1502
rect 13758 1490 13788 1502
rect 13950 1490 13980 1502
rect 14142 1490 14172 1502
rect 14818 1490 14848 1502
rect 15010 1490 15040 1502
rect 15202 1490 15232 1502
rect 15394 1490 15424 1502
rect 15586 1490 15616 1502
rect 15778 1490 15808 1502
rect 15970 1490 16000 1502
rect 16646 1490 16676 1502
rect 16838 1490 16868 1502
rect 17030 1490 17060 1502
rect 17222 1490 17252 1502
rect 17414 1490 17444 1502
rect 17606 1490 17636 1502
rect 17798 1490 17828 1502
rect 18474 1490 18504 1502
rect 18666 1490 18696 1502
rect 18858 1490 18888 1502
rect 19050 1490 19080 1502
rect 19242 1490 19272 1502
rect 19434 1490 19464 1502
rect 19626 1490 19656 1502
rect 20302 1490 20332 1502
rect 20494 1490 20524 1502
rect 20686 1490 20716 1502
rect 20878 1490 20908 1502
rect 21070 1490 21100 1502
rect 21262 1490 21292 1502
rect 21454 1490 21484 1502
rect 0 1431 1490 1490
rect 1828 1431 3318 1490
rect 3656 1431 5146 1490
rect 5484 1431 6974 1490
rect 7312 1431 8802 1490
rect 9140 1431 10630 1490
rect 10968 1431 12458 1490
rect 12796 1431 14286 1490
rect 14624 1431 16114 1490
rect 16452 1431 17942 1490
rect 18280 1431 19770 1490
rect 20108 1431 21598 1490
rect 0 1252 1490 1311
rect 1828 1252 3318 1311
rect 3656 1252 5146 1311
rect 5484 1252 6974 1311
rect 7312 1252 8802 1311
rect 9140 1252 10630 1311
rect 10968 1252 12458 1311
rect 12796 1252 14286 1311
rect 14624 1252 16114 1311
rect 16452 1252 17942 1311
rect 18280 1252 19770 1311
rect 20108 1252 21598 1311
rect 98 1240 128 1252
rect 290 1240 320 1252
rect 482 1240 512 1252
rect 674 1240 704 1252
rect 866 1240 896 1252
rect 1058 1240 1088 1252
rect 1250 1240 1280 1252
rect 1442 1240 1472 1252
rect 1926 1240 1956 1252
rect 2118 1240 2148 1252
rect 2310 1240 2340 1252
rect 2502 1240 2532 1252
rect 2694 1240 2724 1252
rect 2886 1240 2916 1252
rect 3078 1240 3108 1252
rect 3270 1240 3300 1252
rect 3754 1240 3784 1252
rect 3946 1240 3976 1252
rect 4138 1240 4168 1252
rect 4330 1240 4360 1252
rect 4522 1240 4552 1252
rect 4714 1240 4744 1252
rect 4906 1240 4936 1252
rect 5098 1240 5128 1252
rect 5582 1240 5612 1252
rect 5774 1240 5804 1252
rect 5966 1240 5996 1252
rect 6158 1240 6188 1252
rect 6350 1240 6380 1252
rect 6542 1240 6572 1252
rect 6734 1240 6764 1252
rect 6926 1240 6956 1252
rect 7410 1240 7440 1252
rect 7602 1240 7632 1252
rect 7794 1240 7824 1252
rect 7986 1240 8016 1252
rect 8178 1240 8208 1252
rect 8370 1240 8400 1252
rect 8562 1240 8592 1252
rect 8754 1240 8784 1252
rect 9238 1240 9268 1252
rect 9430 1240 9460 1252
rect 9622 1240 9652 1252
rect 9814 1240 9844 1252
rect 10006 1240 10036 1252
rect 10198 1240 10228 1252
rect 10390 1240 10420 1252
rect 10582 1240 10612 1252
rect 11066 1240 11096 1252
rect 11258 1240 11288 1252
rect 11450 1240 11480 1252
rect 11642 1240 11672 1252
rect 11834 1240 11864 1252
rect 12026 1240 12056 1252
rect 12218 1240 12248 1252
rect 12410 1240 12440 1252
rect 12894 1240 12924 1252
rect 13086 1240 13116 1252
rect 13278 1240 13308 1252
rect 13470 1240 13500 1252
rect 13662 1240 13692 1252
rect 13854 1240 13884 1252
rect 14046 1240 14076 1252
rect 14238 1240 14268 1252
rect 14722 1240 14752 1252
rect 14914 1240 14944 1252
rect 15106 1240 15136 1252
rect 15298 1240 15328 1252
rect 15490 1240 15520 1252
rect 15682 1240 15712 1252
rect 15874 1240 15904 1252
rect 16066 1240 16096 1252
rect 16550 1240 16580 1252
rect 16742 1240 16772 1252
rect 16934 1240 16964 1252
rect 17126 1240 17156 1252
rect 17318 1240 17348 1252
rect 17510 1240 17540 1252
rect 17702 1240 17732 1252
rect 17894 1240 17924 1252
rect 18378 1240 18408 1252
rect 18570 1240 18600 1252
rect 18762 1240 18792 1252
rect 18954 1240 18984 1252
rect 19146 1240 19176 1252
rect 19338 1240 19368 1252
rect 19530 1240 19560 1252
rect 19722 1240 19752 1252
rect 20206 1240 20236 1252
rect 20398 1240 20428 1252
rect 20590 1240 20620 1252
rect 20782 1240 20812 1252
rect 20974 1240 21004 1252
rect 21166 1240 21196 1252
rect 21358 1240 21388 1252
rect 21550 1240 21580 1252
rect 194 776 224 788
rect 386 776 416 788
rect 578 776 608 788
rect 770 776 800 788
rect 962 776 992 788
rect 1154 776 1184 788
rect 1346 776 1376 788
rect 2022 776 2052 788
rect 2214 776 2244 788
rect 2406 776 2436 788
rect 2598 776 2628 788
rect 2790 776 2820 788
rect 2982 776 3012 788
rect 3174 776 3204 788
rect 3850 776 3880 788
rect 4042 776 4072 788
rect 4234 776 4264 788
rect 4426 776 4456 788
rect 4618 776 4648 788
rect 4810 776 4840 788
rect 5002 776 5032 788
rect 5678 776 5708 788
rect 5870 776 5900 788
rect 6062 776 6092 788
rect 6254 776 6284 788
rect 6446 776 6476 788
rect 6638 776 6668 788
rect 6830 776 6860 788
rect 7506 776 7536 788
rect 7698 776 7728 788
rect 7890 776 7920 788
rect 8082 776 8112 788
rect 8274 776 8304 788
rect 8466 776 8496 788
rect 8658 776 8688 788
rect 9334 776 9364 788
rect 9526 776 9556 788
rect 9718 776 9748 788
rect 9910 776 9940 788
rect 10102 776 10132 788
rect 10294 776 10324 788
rect 10486 776 10516 788
rect 11162 776 11192 788
rect 11354 776 11384 788
rect 11546 776 11576 788
rect 11738 776 11768 788
rect 11930 776 11960 788
rect 12122 776 12152 788
rect 12314 776 12344 788
rect 12990 776 13020 788
rect 13182 776 13212 788
rect 13374 776 13404 788
rect 13566 776 13596 788
rect 13758 776 13788 788
rect 13950 776 13980 788
rect 14142 776 14172 788
rect 14818 776 14848 788
rect 15010 776 15040 788
rect 15202 776 15232 788
rect 15394 776 15424 788
rect 15586 776 15616 788
rect 15778 776 15808 788
rect 15970 776 16000 788
rect 16646 776 16676 788
rect 16838 776 16868 788
rect 17030 776 17060 788
rect 17222 776 17252 788
rect 17414 776 17444 788
rect 17606 776 17636 788
rect 17798 776 17828 788
rect 18474 776 18504 788
rect 18666 776 18696 788
rect 18858 776 18888 788
rect 19050 776 19080 788
rect 19242 776 19272 788
rect 19434 776 19464 788
rect 19626 776 19656 788
rect 20302 776 20332 788
rect 20494 776 20524 788
rect 20686 776 20716 788
rect 20878 776 20908 788
rect 21070 776 21100 788
rect 21262 776 21292 788
rect 21454 776 21484 788
rect 0 717 1490 776
rect 1828 717 3318 776
rect 3656 717 5146 776
rect 5484 717 6974 776
rect 7312 717 8802 776
rect 9140 717 10630 776
rect 10968 717 12458 776
rect 12796 717 14286 776
rect 14624 717 16114 776
rect 16452 717 17942 776
rect 18280 717 19770 776
rect 20108 717 21598 776
rect 0 538 1490 597
rect 1828 538 3318 597
rect 3656 538 5146 597
rect 5484 538 6974 597
rect 7312 538 8802 597
rect 9140 538 10630 597
rect 10968 538 12458 597
rect 12796 538 14286 597
rect 14624 538 16114 597
rect 16452 538 17942 597
rect 18280 538 19770 597
rect 20108 538 21598 597
rect 98 526 128 538
rect 290 526 320 538
rect 482 526 512 538
rect 674 526 704 538
rect 866 526 896 538
rect 1058 526 1088 538
rect 1250 526 1280 538
rect 1442 526 1472 538
rect 1926 526 1956 538
rect 2118 526 2148 538
rect 2310 526 2340 538
rect 2502 526 2532 538
rect 2694 526 2724 538
rect 2886 526 2916 538
rect 3078 526 3108 538
rect 3270 526 3300 538
rect 3754 526 3784 538
rect 3946 526 3976 538
rect 4138 526 4168 538
rect 4330 526 4360 538
rect 4522 526 4552 538
rect 4714 526 4744 538
rect 4906 526 4936 538
rect 5098 526 5128 538
rect 5582 526 5612 538
rect 5774 526 5804 538
rect 5966 526 5996 538
rect 6158 526 6188 538
rect 6350 526 6380 538
rect 6542 526 6572 538
rect 6734 526 6764 538
rect 6926 526 6956 538
rect 7410 526 7440 538
rect 7602 526 7632 538
rect 7794 526 7824 538
rect 7986 526 8016 538
rect 8178 526 8208 538
rect 8370 526 8400 538
rect 8562 526 8592 538
rect 8754 526 8784 538
rect 9238 526 9268 538
rect 9430 526 9460 538
rect 9622 526 9652 538
rect 9814 526 9844 538
rect 10006 526 10036 538
rect 10198 526 10228 538
rect 10390 526 10420 538
rect 10582 526 10612 538
rect 11066 526 11096 538
rect 11258 526 11288 538
rect 11450 526 11480 538
rect 11642 526 11672 538
rect 11834 526 11864 538
rect 12026 526 12056 538
rect 12218 526 12248 538
rect 12410 526 12440 538
rect 12894 526 12924 538
rect 13086 526 13116 538
rect 13278 526 13308 538
rect 13470 526 13500 538
rect 13662 526 13692 538
rect 13854 526 13884 538
rect 14046 526 14076 538
rect 14238 526 14268 538
rect 14722 526 14752 538
rect 14914 526 14944 538
rect 15106 526 15136 538
rect 15298 526 15328 538
rect 15490 526 15520 538
rect 15682 526 15712 538
rect 15874 526 15904 538
rect 16066 526 16096 538
rect 16550 526 16580 538
rect 16742 526 16772 538
rect 16934 526 16964 538
rect 17126 526 17156 538
rect 17318 526 17348 538
rect 17510 526 17540 538
rect 17702 526 17732 538
rect 17894 526 17924 538
rect 18378 526 18408 538
rect 18570 526 18600 538
rect 18762 526 18792 538
rect 18954 526 18984 538
rect 19146 526 19176 538
rect 19338 526 19368 538
rect 19530 526 19560 538
rect 19722 526 19752 538
rect 20206 526 20236 538
rect 20398 526 20428 538
rect 20590 526 20620 538
rect 20782 526 20812 538
rect 20974 526 21004 538
rect 21166 526 21196 538
rect 21358 526 21388 538
rect 21550 526 21580 538
rect 194 62 224 74
rect 386 62 416 74
rect 578 62 608 74
rect 770 62 800 74
rect 962 62 992 74
rect 1154 62 1184 74
rect 1346 62 1376 74
rect 2022 62 2052 74
rect 2214 62 2244 74
rect 2406 62 2436 74
rect 2598 62 2628 74
rect 2790 62 2820 74
rect 2982 62 3012 74
rect 3174 62 3204 74
rect 3850 62 3880 74
rect 4042 62 4072 74
rect 4234 62 4264 74
rect 4426 62 4456 74
rect 4618 62 4648 74
rect 4810 62 4840 74
rect 5002 62 5032 74
rect 5678 62 5708 74
rect 5870 62 5900 74
rect 6062 62 6092 74
rect 6254 62 6284 74
rect 6446 62 6476 74
rect 6638 62 6668 74
rect 6830 62 6860 74
rect 7506 62 7536 74
rect 7698 62 7728 74
rect 7890 62 7920 74
rect 8082 62 8112 74
rect 8274 62 8304 74
rect 8466 62 8496 74
rect 8658 62 8688 74
rect 9334 62 9364 74
rect 9526 62 9556 74
rect 9718 62 9748 74
rect 9910 62 9940 74
rect 10102 62 10132 74
rect 10294 62 10324 74
rect 10486 62 10516 74
rect 11162 62 11192 74
rect 11354 62 11384 74
rect 11546 62 11576 74
rect 11738 62 11768 74
rect 11930 62 11960 74
rect 12122 62 12152 74
rect 12314 62 12344 74
rect 12990 62 13020 74
rect 13182 62 13212 74
rect 13374 62 13404 74
rect 13566 62 13596 74
rect 13758 62 13788 74
rect 13950 62 13980 74
rect 14142 62 14172 74
rect 14818 62 14848 74
rect 15010 62 15040 74
rect 15202 62 15232 74
rect 15394 62 15424 74
rect 15586 62 15616 74
rect 15778 62 15808 74
rect 15970 62 16000 74
rect 16646 62 16676 74
rect 16838 62 16868 74
rect 17030 62 17060 74
rect 17222 62 17252 74
rect 17414 62 17444 74
rect 17606 62 17636 74
rect 17798 62 17828 74
rect 18474 62 18504 74
rect 18666 62 18696 74
rect 18858 62 18888 74
rect 19050 62 19080 74
rect 19242 62 19272 74
rect 19434 62 19464 74
rect 19626 62 19656 74
rect 20302 62 20332 74
rect 20494 62 20524 74
rect 20686 62 20716 74
rect 20878 62 20908 74
rect 21070 62 21100 74
rect 21262 62 21292 74
rect 21454 62 21484 74
rect 0 3 1490 62
rect 1828 3 3318 62
rect 3656 3 5146 62
rect 5484 3 6974 62
rect 7312 3 8802 62
rect 9140 3 10630 62
rect 10968 3 12458 62
rect 12796 3 14286 62
rect 14624 3 16114 62
rect 16452 3 17942 62
rect 18280 3 19770 62
rect 20108 3 21598 62
<< locali >>
rect 0 21244 1472 21303
rect 1828 21244 3300 21303
rect 3656 21244 5128 21303
rect 5484 21244 6956 21303
rect 7312 21244 8784 21303
rect 9140 21244 10612 21303
rect 10968 21244 12440 21303
rect 12796 21244 14268 21303
rect 14624 21244 16096 21303
rect 16452 21244 17924 21303
rect 18280 21244 19752 21303
rect 20108 21244 21580 21303
rect 1630 21210 1708 21221
rect 3458 21210 3536 21221
rect 5286 21210 5364 21221
rect 7114 21210 7192 21221
rect 8942 21210 9020 21221
rect 10770 21210 10848 21221
rect 12598 21210 12676 21221
rect 14426 21210 14504 21221
rect 16254 21210 16332 21221
rect 18082 21210 18160 21221
rect 19910 21210 19988 21221
rect 21738 21210 21816 21221
rect 1488 21194 1708 21210
rect 1488 20818 1630 21194
rect 1488 20802 1708 20818
rect 3316 21194 3536 21210
rect 3316 20818 3458 21194
rect 3316 20802 3536 20818
rect 5144 21194 5364 21210
rect 5144 20818 5286 21194
rect 5144 20802 5364 20818
rect 6972 21194 7192 21210
rect 6972 20818 7114 21194
rect 6972 20802 7192 20818
rect 8800 21194 9020 21210
rect 8800 20818 8942 21194
rect 8800 20802 9020 20818
rect 10628 21194 10848 21210
rect 10628 20818 10770 21194
rect 10628 20802 10848 20818
rect 12456 21194 12676 21210
rect 12456 20818 12598 21194
rect 12456 20802 12676 20818
rect 14284 21194 14504 21210
rect 14284 20818 14426 21194
rect 14284 20802 14504 20818
rect 16112 21194 16332 21210
rect 16112 20818 16254 21194
rect 16112 20802 16332 20818
rect 17940 21194 18160 21210
rect 17940 20818 18082 21194
rect 17940 20802 18160 20818
rect 19768 21194 19988 21210
rect 19768 20818 19910 21194
rect 19768 20802 19988 20818
rect 21596 21194 21816 21210
rect 21596 20818 21738 21194
rect 21596 20802 21816 20818
rect 1630 20791 1708 20802
rect 3458 20791 3536 20802
rect 5286 20791 5364 20802
rect 7114 20791 7192 20802
rect 8942 20791 9020 20802
rect 10770 20791 10848 20802
rect 12598 20791 12676 20802
rect 14426 20791 14504 20802
rect 16254 20791 16332 20802
rect 18082 20791 18160 20802
rect 19910 20791 19988 20802
rect 21738 20791 21816 20802
rect 0 20709 1490 20768
rect 1828 20709 3318 20768
rect 3656 20709 5146 20768
rect 5484 20709 6974 20768
rect 7312 20709 8802 20768
rect 9140 20709 10630 20768
rect 10968 20709 12458 20768
rect 12796 20709 14286 20768
rect 14624 20709 16114 20768
rect 16452 20709 17942 20768
rect 18280 20709 19770 20768
rect 20108 20709 21598 20768
rect 0 20530 1472 20589
rect 1828 20530 3300 20589
rect 3656 20530 5128 20589
rect 5484 20530 6956 20589
rect 7312 20530 8784 20589
rect 9140 20530 10612 20589
rect 10968 20530 12440 20589
rect 12796 20530 14268 20589
rect 14624 20530 16096 20589
rect 16452 20530 17924 20589
rect 18280 20530 19752 20589
rect 20108 20530 21580 20589
rect 1630 20496 1708 20507
rect 3458 20496 3536 20507
rect 5286 20496 5364 20507
rect 7114 20496 7192 20507
rect 8942 20496 9020 20507
rect 10770 20496 10848 20507
rect 12598 20496 12676 20507
rect 14426 20496 14504 20507
rect 16254 20496 16332 20507
rect 18082 20496 18160 20507
rect 19910 20496 19988 20507
rect 21738 20496 21816 20507
rect 1488 20480 1708 20496
rect 1488 20104 1630 20480
rect 1488 20088 1708 20104
rect 3316 20480 3536 20496
rect 3316 20104 3458 20480
rect 3316 20088 3536 20104
rect 5144 20480 5364 20496
rect 5144 20104 5286 20480
rect 5144 20088 5364 20104
rect 6972 20480 7192 20496
rect 6972 20104 7114 20480
rect 6972 20088 7192 20104
rect 8800 20480 9020 20496
rect 8800 20104 8942 20480
rect 8800 20088 9020 20104
rect 10628 20480 10848 20496
rect 10628 20104 10770 20480
rect 10628 20088 10848 20104
rect 12456 20480 12676 20496
rect 12456 20104 12598 20480
rect 12456 20088 12676 20104
rect 14284 20480 14504 20496
rect 14284 20104 14426 20480
rect 14284 20088 14504 20104
rect 16112 20480 16332 20496
rect 16112 20104 16254 20480
rect 16112 20088 16332 20104
rect 17940 20480 18160 20496
rect 17940 20104 18082 20480
rect 17940 20088 18160 20104
rect 19768 20480 19988 20496
rect 19768 20104 19910 20480
rect 19768 20088 19988 20104
rect 21596 20480 21816 20496
rect 21596 20104 21738 20480
rect 21596 20088 21816 20104
rect 1630 20077 1708 20088
rect 3458 20077 3536 20088
rect 5286 20077 5364 20088
rect 7114 20077 7192 20088
rect 8942 20077 9020 20088
rect 10770 20077 10848 20088
rect 12598 20077 12676 20088
rect 14426 20077 14504 20088
rect 16254 20077 16332 20088
rect 18082 20077 18160 20088
rect 19910 20077 19988 20088
rect 21738 20077 21816 20088
rect 0 19995 1490 20054
rect 1828 19995 3318 20054
rect 3656 19995 5146 20054
rect 5484 19995 6974 20054
rect 7312 19995 8802 20054
rect 9140 19995 10630 20054
rect 10968 19995 12458 20054
rect 12796 19995 14286 20054
rect 14624 19995 16114 20054
rect 16452 19995 17942 20054
rect 18280 19995 19770 20054
rect 20108 19995 21598 20054
rect 0 19816 1472 19875
rect 1828 19816 3300 19875
rect 3656 19816 5128 19875
rect 5484 19816 6956 19875
rect 7312 19816 8784 19875
rect 9140 19816 10612 19875
rect 10968 19816 12440 19875
rect 12796 19816 14268 19875
rect 14624 19816 16096 19875
rect 16452 19816 17924 19875
rect 18280 19816 19752 19875
rect 20108 19816 21580 19875
rect 1630 19782 1708 19793
rect 3458 19782 3536 19793
rect 5286 19782 5364 19793
rect 7114 19782 7192 19793
rect 8942 19782 9020 19793
rect 10770 19782 10848 19793
rect 12598 19782 12676 19793
rect 14426 19782 14504 19793
rect 16254 19782 16332 19793
rect 18082 19782 18160 19793
rect 19910 19782 19988 19793
rect 21738 19782 21816 19793
rect 1488 19766 1708 19782
rect 1488 19390 1630 19766
rect 1488 19374 1708 19390
rect 3316 19766 3536 19782
rect 3316 19390 3458 19766
rect 3316 19374 3536 19390
rect 5144 19766 5364 19782
rect 5144 19390 5286 19766
rect 5144 19374 5364 19390
rect 6972 19766 7192 19782
rect 6972 19390 7114 19766
rect 6972 19374 7192 19390
rect 8800 19766 9020 19782
rect 8800 19390 8942 19766
rect 8800 19374 9020 19390
rect 10628 19766 10848 19782
rect 10628 19390 10770 19766
rect 10628 19374 10848 19390
rect 12456 19766 12676 19782
rect 12456 19390 12598 19766
rect 12456 19374 12676 19390
rect 14284 19766 14504 19782
rect 14284 19390 14426 19766
rect 14284 19374 14504 19390
rect 16112 19766 16332 19782
rect 16112 19390 16254 19766
rect 16112 19374 16332 19390
rect 17940 19766 18160 19782
rect 17940 19390 18082 19766
rect 17940 19374 18160 19390
rect 19768 19766 19988 19782
rect 19768 19390 19910 19766
rect 19768 19374 19988 19390
rect 21596 19766 21816 19782
rect 21596 19390 21738 19766
rect 21596 19374 21816 19390
rect 1630 19363 1708 19374
rect 3458 19363 3536 19374
rect 5286 19363 5364 19374
rect 7114 19363 7192 19374
rect 8942 19363 9020 19374
rect 10770 19363 10848 19374
rect 12598 19363 12676 19374
rect 14426 19363 14504 19374
rect 16254 19363 16332 19374
rect 18082 19363 18160 19374
rect 19910 19363 19988 19374
rect 21738 19363 21816 19374
rect 0 19281 1490 19340
rect 1828 19281 3318 19340
rect 3656 19281 5146 19340
rect 5484 19281 6974 19340
rect 7312 19281 8802 19340
rect 9140 19281 10630 19340
rect 10968 19281 12458 19340
rect 12796 19281 14286 19340
rect 14624 19281 16114 19340
rect 16452 19281 17942 19340
rect 18280 19281 19770 19340
rect 20108 19281 21598 19340
rect 0 19102 1472 19161
rect 1828 19102 3300 19161
rect 3656 19102 5128 19161
rect 5484 19102 6956 19161
rect 7312 19102 8784 19161
rect 9140 19102 10612 19161
rect 10968 19102 12440 19161
rect 12796 19102 14268 19161
rect 14624 19102 16096 19161
rect 16452 19102 17924 19161
rect 18280 19102 19752 19161
rect 20108 19102 21580 19161
rect 1630 19068 1708 19079
rect 3458 19068 3536 19079
rect 5286 19068 5364 19079
rect 7114 19068 7192 19079
rect 8942 19068 9020 19079
rect 10770 19068 10848 19079
rect 12598 19068 12676 19079
rect 14426 19068 14504 19079
rect 16254 19068 16332 19079
rect 18082 19068 18160 19079
rect 19910 19068 19988 19079
rect 21738 19068 21816 19079
rect 1488 19052 1708 19068
rect 1488 18676 1630 19052
rect 1488 18660 1708 18676
rect 3316 19052 3536 19068
rect 3316 18676 3458 19052
rect 3316 18660 3536 18676
rect 5144 19052 5364 19068
rect 5144 18676 5286 19052
rect 5144 18660 5364 18676
rect 6972 19052 7192 19068
rect 6972 18676 7114 19052
rect 6972 18660 7192 18676
rect 8800 19052 9020 19068
rect 8800 18676 8942 19052
rect 8800 18660 9020 18676
rect 10628 19052 10848 19068
rect 10628 18676 10770 19052
rect 10628 18660 10848 18676
rect 12456 19052 12676 19068
rect 12456 18676 12598 19052
rect 12456 18660 12676 18676
rect 14284 19052 14504 19068
rect 14284 18676 14426 19052
rect 14284 18660 14504 18676
rect 16112 19052 16332 19068
rect 16112 18676 16254 19052
rect 16112 18660 16332 18676
rect 17940 19052 18160 19068
rect 17940 18676 18082 19052
rect 17940 18660 18160 18676
rect 19768 19052 19988 19068
rect 19768 18676 19910 19052
rect 19768 18660 19988 18676
rect 21596 19052 21816 19068
rect 21596 18676 21738 19052
rect 21596 18660 21816 18676
rect 1630 18649 1708 18660
rect 3458 18649 3536 18660
rect 5286 18649 5364 18660
rect 7114 18649 7192 18660
rect 8942 18649 9020 18660
rect 10770 18649 10848 18660
rect 12598 18649 12676 18660
rect 14426 18649 14504 18660
rect 16254 18649 16332 18660
rect 18082 18649 18160 18660
rect 19910 18649 19988 18660
rect 21738 18649 21816 18660
rect 0 18567 1490 18626
rect 1828 18567 3318 18626
rect 3656 18567 5146 18626
rect 5484 18567 6974 18626
rect 7312 18567 8802 18626
rect 9140 18567 10630 18626
rect 10968 18567 12458 18626
rect 12796 18567 14286 18626
rect 14624 18567 16114 18626
rect 16452 18567 17942 18626
rect 18280 18567 19770 18626
rect 20108 18567 21598 18626
rect 0 18388 1472 18447
rect 1828 18388 3300 18447
rect 3656 18388 5128 18447
rect 5484 18388 6956 18447
rect 7312 18388 8784 18447
rect 9140 18388 10612 18447
rect 10968 18388 12440 18447
rect 12796 18388 14268 18447
rect 14624 18388 16096 18447
rect 16452 18388 17924 18447
rect 18280 18388 19752 18447
rect 20108 18388 21580 18447
rect 1630 18354 1708 18365
rect 3458 18354 3536 18365
rect 5286 18354 5364 18365
rect 7114 18354 7192 18365
rect 8942 18354 9020 18365
rect 10770 18354 10848 18365
rect 12598 18354 12676 18365
rect 14426 18354 14504 18365
rect 16254 18354 16332 18365
rect 18082 18354 18160 18365
rect 19910 18354 19988 18365
rect 21738 18354 21816 18365
rect 1488 18338 1708 18354
rect 1488 17962 1630 18338
rect 1488 17946 1708 17962
rect 3316 18338 3536 18354
rect 3316 17962 3458 18338
rect 3316 17946 3536 17962
rect 5144 18338 5364 18354
rect 5144 17962 5286 18338
rect 5144 17946 5364 17962
rect 6972 18338 7192 18354
rect 6972 17962 7114 18338
rect 6972 17946 7192 17962
rect 8800 18338 9020 18354
rect 8800 17962 8942 18338
rect 8800 17946 9020 17962
rect 10628 18338 10848 18354
rect 10628 17962 10770 18338
rect 10628 17946 10848 17962
rect 12456 18338 12676 18354
rect 12456 17962 12598 18338
rect 12456 17946 12676 17962
rect 14284 18338 14504 18354
rect 14284 17962 14426 18338
rect 14284 17946 14504 17962
rect 16112 18338 16332 18354
rect 16112 17962 16254 18338
rect 16112 17946 16332 17962
rect 17940 18338 18160 18354
rect 17940 17962 18082 18338
rect 17940 17946 18160 17962
rect 19768 18338 19988 18354
rect 19768 17962 19910 18338
rect 19768 17946 19988 17962
rect 21596 18338 21816 18354
rect 21596 17962 21738 18338
rect 21596 17946 21816 17962
rect 1630 17935 1708 17946
rect 3458 17935 3536 17946
rect 5286 17935 5364 17946
rect 7114 17935 7192 17946
rect 8942 17935 9020 17946
rect 10770 17935 10848 17946
rect 12598 17935 12676 17946
rect 14426 17935 14504 17946
rect 16254 17935 16332 17946
rect 18082 17935 18160 17946
rect 19910 17935 19988 17946
rect 21738 17935 21816 17946
rect 0 17853 1490 17912
rect 1828 17853 3318 17912
rect 3656 17853 5146 17912
rect 5484 17853 6974 17912
rect 7312 17853 8802 17912
rect 9140 17853 10630 17912
rect 10968 17853 12458 17912
rect 12796 17853 14286 17912
rect 14624 17853 16114 17912
rect 16452 17853 17942 17912
rect 18280 17853 19770 17912
rect 20108 17853 21598 17912
rect 0 17674 1472 17733
rect 1828 17674 3300 17733
rect 3656 17674 5128 17733
rect 5484 17674 6956 17733
rect 7312 17674 8784 17733
rect 9140 17674 10612 17733
rect 10968 17674 12440 17733
rect 12796 17674 14268 17733
rect 14624 17674 16096 17733
rect 16452 17674 17924 17733
rect 18280 17674 19752 17733
rect 20108 17674 21580 17733
rect 1630 17640 1708 17651
rect 3458 17640 3536 17651
rect 5286 17640 5364 17651
rect 7114 17640 7192 17651
rect 8942 17640 9020 17651
rect 10770 17640 10848 17651
rect 12598 17640 12676 17651
rect 14426 17640 14504 17651
rect 16254 17640 16332 17651
rect 18082 17640 18160 17651
rect 19910 17640 19988 17651
rect 21738 17640 21816 17651
rect 1488 17624 1708 17640
rect 1488 17248 1630 17624
rect 1488 17232 1708 17248
rect 3316 17624 3536 17640
rect 3316 17248 3458 17624
rect 3316 17232 3536 17248
rect 5144 17624 5364 17640
rect 5144 17248 5286 17624
rect 5144 17232 5364 17248
rect 6972 17624 7192 17640
rect 6972 17248 7114 17624
rect 6972 17232 7192 17248
rect 8800 17624 9020 17640
rect 8800 17248 8942 17624
rect 8800 17232 9020 17248
rect 10628 17624 10848 17640
rect 10628 17248 10770 17624
rect 10628 17232 10848 17248
rect 12456 17624 12676 17640
rect 12456 17248 12598 17624
rect 12456 17232 12676 17248
rect 14284 17624 14504 17640
rect 14284 17248 14426 17624
rect 14284 17232 14504 17248
rect 16112 17624 16332 17640
rect 16112 17248 16254 17624
rect 16112 17232 16332 17248
rect 17940 17624 18160 17640
rect 17940 17248 18082 17624
rect 17940 17232 18160 17248
rect 19768 17624 19988 17640
rect 19768 17248 19910 17624
rect 19768 17232 19988 17248
rect 21596 17624 21816 17640
rect 21596 17248 21738 17624
rect 21596 17232 21816 17248
rect 1630 17221 1708 17232
rect 3458 17221 3536 17232
rect 5286 17221 5364 17232
rect 7114 17221 7192 17232
rect 8942 17221 9020 17232
rect 10770 17221 10848 17232
rect 12598 17221 12676 17232
rect 14426 17221 14504 17232
rect 16254 17221 16332 17232
rect 18082 17221 18160 17232
rect 19910 17221 19988 17232
rect 21738 17221 21816 17232
rect 0 17139 1490 17198
rect 1828 17139 3318 17198
rect 3656 17139 5146 17198
rect 5484 17139 6974 17198
rect 7312 17139 8802 17198
rect 9140 17139 10630 17198
rect 10968 17139 12458 17198
rect 12796 17139 14286 17198
rect 14624 17139 16114 17198
rect 16452 17139 17942 17198
rect 18280 17139 19770 17198
rect 20108 17139 21598 17198
rect 0 16960 1472 17019
rect 1828 16960 3300 17019
rect 3656 16960 5128 17019
rect 5484 16960 6956 17019
rect 7312 16960 8784 17019
rect 9140 16960 10612 17019
rect 10968 16960 12440 17019
rect 12796 16960 14268 17019
rect 14624 16960 16096 17019
rect 16452 16960 17924 17019
rect 18280 16960 19752 17019
rect 20108 16960 21580 17019
rect 1630 16926 1708 16937
rect 3458 16926 3536 16937
rect 5286 16926 5364 16937
rect 7114 16926 7192 16937
rect 8942 16926 9020 16937
rect 10770 16926 10848 16937
rect 12598 16926 12676 16937
rect 14426 16926 14504 16937
rect 16254 16926 16332 16937
rect 18082 16926 18160 16937
rect 19910 16926 19988 16937
rect 21738 16926 21816 16937
rect 1488 16910 1708 16926
rect 1488 16534 1630 16910
rect 1488 16518 1708 16534
rect 3316 16910 3536 16926
rect 3316 16534 3458 16910
rect 3316 16518 3536 16534
rect 5144 16910 5364 16926
rect 5144 16534 5286 16910
rect 5144 16518 5364 16534
rect 6972 16910 7192 16926
rect 6972 16534 7114 16910
rect 6972 16518 7192 16534
rect 8800 16910 9020 16926
rect 8800 16534 8942 16910
rect 8800 16518 9020 16534
rect 10628 16910 10848 16926
rect 10628 16534 10770 16910
rect 10628 16518 10848 16534
rect 12456 16910 12676 16926
rect 12456 16534 12598 16910
rect 12456 16518 12676 16534
rect 14284 16910 14504 16926
rect 14284 16534 14426 16910
rect 14284 16518 14504 16534
rect 16112 16910 16332 16926
rect 16112 16534 16254 16910
rect 16112 16518 16332 16534
rect 17940 16910 18160 16926
rect 17940 16534 18082 16910
rect 17940 16518 18160 16534
rect 19768 16910 19988 16926
rect 19768 16534 19910 16910
rect 19768 16518 19988 16534
rect 21596 16910 21816 16926
rect 21596 16534 21738 16910
rect 21596 16518 21816 16534
rect 1630 16507 1708 16518
rect 3458 16507 3536 16518
rect 5286 16507 5364 16518
rect 7114 16507 7192 16518
rect 8942 16507 9020 16518
rect 10770 16507 10848 16518
rect 12598 16507 12676 16518
rect 14426 16507 14504 16518
rect 16254 16507 16332 16518
rect 18082 16507 18160 16518
rect 19910 16507 19988 16518
rect 21738 16507 21816 16518
rect 0 16425 1490 16484
rect 1828 16425 3318 16484
rect 3656 16425 5146 16484
rect 5484 16425 6974 16484
rect 7312 16425 8802 16484
rect 9140 16425 10630 16484
rect 10968 16425 12458 16484
rect 12796 16425 14286 16484
rect 14624 16425 16114 16484
rect 16452 16425 17942 16484
rect 18280 16425 19770 16484
rect 20108 16425 21598 16484
rect 0 16246 1472 16305
rect 1828 16246 3300 16305
rect 3656 16246 5128 16305
rect 5484 16246 6956 16305
rect 7312 16246 8784 16305
rect 9140 16246 10612 16305
rect 10968 16246 12440 16305
rect 12796 16246 14268 16305
rect 14624 16246 16096 16305
rect 16452 16246 17924 16305
rect 18280 16246 19752 16305
rect 20108 16246 21580 16305
rect 1630 16212 1708 16223
rect 3458 16212 3536 16223
rect 5286 16212 5364 16223
rect 7114 16212 7192 16223
rect 8942 16212 9020 16223
rect 10770 16212 10848 16223
rect 12598 16212 12676 16223
rect 14426 16212 14504 16223
rect 16254 16212 16332 16223
rect 18082 16212 18160 16223
rect 19910 16212 19988 16223
rect 21738 16212 21816 16223
rect 1488 16196 1708 16212
rect 1488 15820 1630 16196
rect 1488 15804 1708 15820
rect 3316 16196 3536 16212
rect 3316 15820 3458 16196
rect 3316 15804 3536 15820
rect 5144 16196 5364 16212
rect 5144 15820 5286 16196
rect 5144 15804 5364 15820
rect 6972 16196 7192 16212
rect 6972 15820 7114 16196
rect 6972 15804 7192 15820
rect 8800 16196 9020 16212
rect 8800 15820 8942 16196
rect 8800 15804 9020 15820
rect 10628 16196 10848 16212
rect 10628 15820 10770 16196
rect 10628 15804 10848 15820
rect 12456 16196 12676 16212
rect 12456 15820 12598 16196
rect 12456 15804 12676 15820
rect 14284 16196 14504 16212
rect 14284 15820 14426 16196
rect 14284 15804 14504 15820
rect 16112 16196 16332 16212
rect 16112 15820 16254 16196
rect 16112 15804 16332 15820
rect 17940 16196 18160 16212
rect 17940 15820 18082 16196
rect 17940 15804 18160 15820
rect 19768 16196 19988 16212
rect 19768 15820 19910 16196
rect 19768 15804 19988 15820
rect 21596 16196 21816 16212
rect 21596 15820 21738 16196
rect 21596 15804 21816 15820
rect 1630 15793 1708 15804
rect 3458 15793 3536 15804
rect 5286 15793 5364 15804
rect 7114 15793 7192 15804
rect 8942 15793 9020 15804
rect 10770 15793 10848 15804
rect 12598 15793 12676 15804
rect 14426 15793 14504 15804
rect 16254 15793 16332 15804
rect 18082 15793 18160 15804
rect 19910 15793 19988 15804
rect 21738 15793 21816 15804
rect 0 15711 1490 15770
rect 1828 15711 3318 15770
rect 3656 15711 5146 15770
rect 5484 15711 6974 15770
rect 7312 15711 8802 15770
rect 9140 15711 10630 15770
rect 10968 15711 12458 15770
rect 12796 15711 14286 15770
rect 14624 15711 16114 15770
rect 16452 15711 17942 15770
rect 18280 15711 19770 15770
rect 20108 15711 21598 15770
rect 0 15532 1472 15591
rect 1828 15532 3300 15591
rect 3656 15532 5128 15591
rect 5484 15532 6956 15591
rect 7312 15532 8784 15591
rect 9140 15532 10612 15591
rect 10968 15532 12440 15591
rect 12796 15532 14268 15591
rect 14624 15532 16096 15591
rect 16452 15532 17924 15591
rect 18280 15532 19752 15591
rect 20108 15532 21580 15591
rect 1630 15498 1708 15509
rect 3458 15498 3536 15509
rect 5286 15498 5364 15509
rect 7114 15498 7192 15509
rect 8942 15498 9020 15509
rect 10770 15498 10848 15509
rect 12598 15498 12676 15509
rect 14426 15498 14504 15509
rect 16254 15498 16332 15509
rect 18082 15498 18160 15509
rect 19910 15498 19988 15509
rect 21738 15498 21816 15509
rect 1488 15482 1708 15498
rect 1488 15106 1630 15482
rect 1488 15090 1708 15106
rect 3316 15482 3536 15498
rect 3316 15106 3458 15482
rect 3316 15090 3536 15106
rect 5144 15482 5364 15498
rect 5144 15106 5286 15482
rect 5144 15090 5364 15106
rect 6972 15482 7192 15498
rect 6972 15106 7114 15482
rect 6972 15090 7192 15106
rect 8800 15482 9020 15498
rect 8800 15106 8942 15482
rect 8800 15090 9020 15106
rect 10628 15482 10848 15498
rect 10628 15106 10770 15482
rect 10628 15090 10848 15106
rect 12456 15482 12676 15498
rect 12456 15106 12598 15482
rect 12456 15090 12676 15106
rect 14284 15482 14504 15498
rect 14284 15106 14426 15482
rect 14284 15090 14504 15106
rect 16112 15482 16332 15498
rect 16112 15106 16254 15482
rect 16112 15090 16332 15106
rect 17940 15482 18160 15498
rect 17940 15106 18082 15482
rect 17940 15090 18160 15106
rect 19768 15482 19988 15498
rect 19768 15106 19910 15482
rect 19768 15090 19988 15106
rect 21596 15482 21816 15498
rect 21596 15106 21738 15482
rect 21596 15090 21816 15106
rect 1630 15079 1708 15090
rect 3458 15079 3536 15090
rect 5286 15079 5364 15090
rect 7114 15079 7192 15090
rect 8942 15079 9020 15090
rect 10770 15079 10848 15090
rect 12598 15079 12676 15090
rect 14426 15079 14504 15090
rect 16254 15079 16332 15090
rect 18082 15079 18160 15090
rect 19910 15079 19988 15090
rect 21738 15079 21816 15090
rect 0 14997 1490 15056
rect 1828 14997 3318 15056
rect 3656 14997 5146 15056
rect 5484 14997 6974 15056
rect 7312 14997 8802 15056
rect 9140 14997 10630 15056
rect 10968 14997 12458 15056
rect 12796 14997 14286 15056
rect 14624 14997 16114 15056
rect 16452 14997 17942 15056
rect 18280 14997 19770 15056
rect 20108 14997 21598 15056
rect 0 14818 1472 14877
rect 1828 14818 3300 14877
rect 3656 14818 5128 14877
rect 5484 14818 6956 14877
rect 7312 14818 8784 14877
rect 9140 14818 10612 14877
rect 10968 14818 12440 14877
rect 12796 14818 14268 14877
rect 14624 14818 16096 14877
rect 16452 14818 17924 14877
rect 18280 14818 19752 14877
rect 20108 14818 21580 14877
rect 1630 14784 1708 14795
rect 3458 14784 3536 14795
rect 5286 14784 5364 14795
rect 7114 14784 7192 14795
rect 8942 14784 9020 14795
rect 10770 14784 10848 14795
rect 12598 14784 12676 14795
rect 14426 14784 14504 14795
rect 16254 14784 16332 14795
rect 18082 14784 18160 14795
rect 19910 14784 19988 14795
rect 21738 14784 21816 14795
rect 1488 14768 1708 14784
rect 1488 14392 1630 14768
rect 1488 14376 1708 14392
rect 3316 14768 3536 14784
rect 3316 14392 3458 14768
rect 3316 14376 3536 14392
rect 5144 14768 5364 14784
rect 5144 14392 5286 14768
rect 5144 14376 5364 14392
rect 6972 14768 7192 14784
rect 6972 14392 7114 14768
rect 6972 14376 7192 14392
rect 8800 14768 9020 14784
rect 8800 14392 8942 14768
rect 8800 14376 9020 14392
rect 10628 14768 10848 14784
rect 10628 14392 10770 14768
rect 10628 14376 10848 14392
rect 12456 14768 12676 14784
rect 12456 14392 12598 14768
rect 12456 14376 12676 14392
rect 14284 14768 14504 14784
rect 14284 14392 14426 14768
rect 14284 14376 14504 14392
rect 16112 14768 16332 14784
rect 16112 14392 16254 14768
rect 16112 14376 16332 14392
rect 17940 14768 18160 14784
rect 17940 14392 18082 14768
rect 17940 14376 18160 14392
rect 19768 14768 19988 14784
rect 19768 14392 19910 14768
rect 19768 14376 19988 14392
rect 21596 14768 21816 14784
rect 21596 14392 21738 14768
rect 21596 14376 21816 14392
rect 1630 14365 1708 14376
rect 3458 14365 3536 14376
rect 5286 14365 5364 14376
rect 7114 14365 7192 14376
rect 8942 14365 9020 14376
rect 10770 14365 10848 14376
rect 12598 14365 12676 14376
rect 14426 14365 14504 14376
rect 16254 14365 16332 14376
rect 18082 14365 18160 14376
rect 19910 14365 19988 14376
rect 21738 14365 21816 14376
rect 0 14283 1490 14342
rect 1828 14283 3318 14342
rect 3656 14283 5146 14342
rect 5484 14283 6974 14342
rect 7312 14283 8802 14342
rect 9140 14283 10630 14342
rect 10968 14283 12458 14342
rect 12796 14283 14286 14342
rect 14624 14283 16114 14342
rect 16452 14283 17942 14342
rect 18280 14283 19770 14342
rect 20108 14283 21598 14342
rect 0 14104 1472 14163
rect 1828 14104 3300 14163
rect 3656 14104 5128 14163
rect 5484 14104 6956 14163
rect 7312 14104 8784 14163
rect 9140 14104 10612 14163
rect 10968 14104 12440 14163
rect 12796 14104 14268 14163
rect 14624 14104 16096 14163
rect 16452 14104 17924 14163
rect 18280 14104 19752 14163
rect 20108 14104 21580 14163
rect 1630 14070 1708 14081
rect 3458 14070 3536 14081
rect 5286 14070 5364 14081
rect 7114 14070 7192 14081
rect 8942 14070 9020 14081
rect 10770 14070 10848 14081
rect 12598 14070 12676 14081
rect 14426 14070 14504 14081
rect 16254 14070 16332 14081
rect 18082 14070 18160 14081
rect 19910 14070 19988 14081
rect 21738 14070 21816 14081
rect 1488 14054 1708 14070
rect 1488 13678 1630 14054
rect 1488 13662 1708 13678
rect 3316 14054 3536 14070
rect 3316 13678 3458 14054
rect 3316 13662 3536 13678
rect 5144 14054 5364 14070
rect 5144 13678 5286 14054
rect 5144 13662 5364 13678
rect 6972 14054 7192 14070
rect 6972 13678 7114 14054
rect 6972 13662 7192 13678
rect 8800 14054 9020 14070
rect 8800 13678 8942 14054
rect 8800 13662 9020 13678
rect 10628 14054 10848 14070
rect 10628 13678 10770 14054
rect 10628 13662 10848 13678
rect 12456 14054 12676 14070
rect 12456 13678 12598 14054
rect 12456 13662 12676 13678
rect 14284 14054 14504 14070
rect 14284 13678 14426 14054
rect 14284 13662 14504 13678
rect 16112 14054 16332 14070
rect 16112 13678 16254 14054
rect 16112 13662 16332 13678
rect 17940 14054 18160 14070
rect 17940 13678 18082 14054
rect 17940 13662 18160 13678
rect 19768 14054 19988 14070
rect 19768 13678 19910 14054
rect 19768 13662 19988 13678
rect 21596 14054 21816 14070
rect 21596 13678 21738 14054
rect 21596 13662 21816 13678
rect 1630 13651 1708 13662
rect 3458 13651 3536 13662
rect 5286 13651 5364 13662
rect 7114 13651 7192 13662
rect 8942 13651 9020 13662
rect 10770 13651 10848 13662
rect 12598 13651 12676 13662
rect 14426 13651 14504 13662
rect 16254 13651 16332 13662
rect 18082 13651 18160 13662
rect 19910 13651 19988 13662
rect 21738 13651 21816 13662
rect 0 13569 1490 13628
rect 1828 13569 3318 13628
rect 3656 13569 5146 13628
rect 5484 13569 6974 13628
rect 7312 13569 8802 13628
rect 9140 13569 10630 13628
rect 10968 13569 12458 13628
rect 12796 13569 14286 13628
rect 14624 13569 16114 13628
rect 16452 13569 17942 13628
rect 18280 13569 19770 13628
rect 20108 13569 21598 13628
rect 0 13390 1472 13449
rect 1828 13390 3300 13449
rect 3656 13390 5128 13449
rect 5484 13390 6956 13449
rect 7312 13390 8784 13449
rect 9140 13390 10612 13449
rect 10968 13390 12440 13449
rect 12796 13390 14268 13449
rect 14624 13390 16096 13449
rect 16452 13390 17924 13449
rect 18280 13390 19752 13449
rect 20108 13390 21580 13449
rect 1630 13356 1708 13367
rect 3458 13356 3536 13367
rect 5286 13356 5364 13367
rect 7114 13356 7192 13367
rect 8942 13356 9020 13367
rect 10770 13356 10848 13367
rect 12598 13356 12676 13367
rect 14426 13356 14504 13367
rect 16254 13356 16332 13367
rect 18082 13356 18160 13367
rect 19910 13356 19988 13367
rect 21738 13356 21816 13367
rect 1488 13340 1708 13356
rect 1488 12964 1630 13340
rect 1488 12948 1708 12964
rect 3316 13340 3536 13356
rect 3316 12964 3458 13340
rect 3316 12948 3536 12964
rect 5144 13340 5364 13356
rect 5144 12964 5286 13340
rect 5144 12948 5364 12964
rect 6972 13340 7192 13356
rect 6972 12964 7114 13340
rect 6972 12948 7192 12964
rect 8800 13340 9020 13356
rect 8800 12964 8942 13340
rect 8800 12948 9020 12964
rect 10628 13340 10848 13356
rect 10628 12964 10770 13340
rect 10628 12948 10848 12964
rect 12456 13340 12676 13356
rect 12456 12964 12598 13340
rect 12456 12948 12676 12964
rect 14284 13340 14504 13356
rect 14284 12964 14426 13340
rect 14284 12948 14504 12964
rect 16112 13340 16332 13356
rect 16112 12964 16254 13340
rect 16112 12948 16332 12964
rect 17940 13340 18160 13356
rect 17940 12964 18082 13340
rect 17940 12948 18160 12964
rect 19768 13340 19988 13356
rect 19768 12964 19910 13340
rect 19768 12948 19988 12964
rect 21596 13340 21816 13356
rect 21596 12964 21738 13340
rect 21596 12948 21816 12964
rect 1630 12937 1708 12948
rect 3458 12937 3536 12948
rect 5286 12937 5364 12948
rect 7114 12937 7192 12948
rect 8942 12937 9020 12948
rect 10770 12937 10848 12948
rect 12598 12937 12676 12948
rect 14426 12937 14504 12948
rect 16254 12937 16332 12948
rect 18082 12937 18160 12948
rect 19910 12937 19988 12948
rect 21738 12937 21816 12948
rect 0 12855 1490 12914
rect 1828 12855 3318 12914
rect 3656 12855 5146 12914
rect 5484 12855 6974 12914
rect 7312 12855 8802 12914
rect 9140 12855 10630 12914
rect 10968 12855 12458 12914
rect 12796 12855 14286 12914
rect 14624 12855 16114 12914
rect 16452 12855 17942 12914
rect 18280 12855 19770 12914
rect 20108 12855 21598 12914
rect 0 12676 1472 12735
rect 1828 12676 3300 12735
rect 3656 12676 5128 12735
rect 5484 12676 6956 12735
rect 7312 12676 8784 12735
rect 9140 12676 10612 12735
rect 10968 12676 12440 12735
rect 12796 12676 14268 12735
rect 14624 12676 16096 12735
rect 16452 12676 17924 12735
rect 18280 12676 19752 12735
rect 20108 12676 21580 12735
rect 1630 12642 1708 12653
rect 3458 12642 3536 12653
rect 5286 12642 5364 12653
rect 7114 12642 7192 12653
rect 8942 12642 9020 12653
rect 10770 12642 10848 12653
rect 12598 12642 12676 12653
rect 14426 12642 14504 12653
rect 16254 12642 16332 12653
rect 18082 12642 18160 12653
rect 19910 12642 19988 12653
rect 21738 12642 21816 12653
rect 1488 12626 1708 12642
rect 1488 12250 1630 12626
rect 1488 12234 1708 12250
rect 3316 12626 3536 12642
rect 3316 12250 3458 12626
rect 3316 12234 3536 12250
rect 5144 12626 5364 12642
rect 5144 12250 5286 12626
rect 5144 12234 5364 12250
rect 6972 12626 7192 12642
rect 6972 12250 7114 12626
rect 6972 12234 7192 12250
rect 8800 12626 9020 12642
rect 8800 12250 8942 12626
rect 8800 12234 9020 12250
rect 10628 12626 10848 12642
rect 10628 12250 10770 12626
rect 10628 12234 10848 12250
rect 12456 12626 12676 12642
rect 12456 12250 12598 12626
rect 12456 12234 12676 12250
rect 14284 12626 14504 12642
rect 14284 12250 14426 12626
rect 14284 12234 14504 12250
rect 16112 12626 16332 12642
rect 16112 12250 16254 12626
rect 16112 12234 16332 12250
rect 17940 12626 18160 12642
rect 17940 12250 18082 12626
rect 17940 12234 18160 12250
rect 19768 12626 19988 12642
rect 19768 12250 19910 12626
rect 19768 12234 19988 12250
rect 21596 12626 21816 12642
rect 21596 12250 21738 12626
rect 21596 12234 21816 12250
rect 1630 12223 1708 12234
rect 3458 12223 3536 12234
rect 5286 12223 5364 12234
rect 7114 12223 7192 12234
rect 8942 12223 9020 12234
rect 10770 12223 10848 12234
rect 12598 12223 12676 12234
rect 14426 12223 14504 12234
rect 16254 12223 16332 12234
rect 18082 12223 18160 12234
rect 19910 12223 19988 12234
rect 21738 12223 21816 12234
rect 0 12141 1490 12200
rect 1828 12141 3318 12200
rect 3656 12141 5146 12200
rect 5484 12141 6974 12200
rect 7312 12141 8802 12200
rect 9140 12141 10630 12200
rect 10968 12141 12458 12200
rect 12796 12141 14286 12200
rect 14624 12141 16114 12200
rect 16452 12141 17942 12200
rect 18280 12141 19770 12200
rect 20108 12141 21598 12200
rect 0 11962 1472 12021
rect 1828 11962 3300 12021
rect 3656 11962 5128 12021
rect 5484 11962 6956 12021
rect 7312 11962 8784 12021
rect 9140 11962 10612 12021
rect 10968 11962 12440 12021
rect 12796 11962 14268 12021
rect 14624 11962 16096 12021
rect 16452 11962 17924 12021
rect 18280 11962 19752 12021
rect 20108 11962 21580 12021
rect 1630 11928 1708 11939
rect 3458 11928 3536 11939
rect 5286 11928 5364 11939
rect 7114 11928 7192 11939
rect 8942 11928 9020 11939
rect 10770 11928 10848 11939
rect 12598 11928 12676 11939
rect 14426 11928 14504 11939
rect 16254 11928 16332 11939
rect 18082 11928 18160 11939
rect 19910 11928 19988 11939
rect 21738 11928 21816 11939
rect 1488 11912 1708 11928
rect 1488 11536 1630 11912
rect 1488 11520 1708 11536
rect 3316 11912 3536 11928
rect 3316 11536 3458 11912
rect 3316 11520 3536 11536
rect 5144 11912 5364 11928
rect 5144 11536 5286 11912
rect 5144 11520 5364 11536
rect 6972 11912 7192 11928
rect 6972 11536 7114 11912
rect 6972 11520 7192 11536
rect 8800 11912 9020 11928
rect 8800 11536 8942 11912
rect 8800 11520 9020 11536
rect 10628 11912 10848 11928
rect 10628 11536 10770 11912
rect 10628 11520 10848 11536
rect 12456 11912 12676 11928
rect 12456 11536 12598 11912
rect 12456 11520 12676 11536
rect 14284 11912 14504 11928
rect 14284 11536 14426 11912
rect 14284 11520 14504 11536
rect 16112 11912 16332 11928
rect 16112 11536 16254 11912
rect 16112 11520 16332 11536
rect 17940 11912 18160 11928
rect 17940 11536 18082 11912
rect 17940 11520 18160 11536
rect 19768 11912 19988 11928
rect 19768 11536 19910 11912
rect 19768 11520 19988 11536
rect 21596 11912 21816 11928
rect 21596 11536 21738 11912
rect 21596 11520 21816 11536
rect 1630 11509 1708 11520
rect 3458 11509 3536 11520
rect 5286 11509 5364 11520
rect 7114 11509 7192 11520
rect 8942 11509 9020 11520
rect 10770 11509 10848 11520
rect 12598 11509 12676 11520
rect 14426 11509 14504 11520
rect 16254 11509 16332 11520
rect 18082 11509 18160 11520
rect 19910 11509 19988 11520
rect 21738 11509 21816 11520
rect 0 11427 1490 11486
rect 1828 11427 3318 11486
rect 3656 11427 5146 11486
rect 5484 11427 6974 11486
rect 7312 11427 8802 11486
rect 9140 11427 10630 11486
rect 10968 11427 12458 11486
rect 12796 11427 14286 11486
rect 14624 11427 16114 11486
rect 16452 11427 17942 11486
rect 18280 11427 19770 11486
rect 20108 11427 21598 11486
rect 0 11248 1472 11307
rect 1828 11248 3300 11307
rect 3656 11248 5128 11307
rect 5484 11248 6956 11307
rect 7312 11248 8784 11307
rect 9140 11248 10612 11307
rect 10968 11248 12440 11307
rect 12796 11248 14268 11307
rect 14624 11248 16096 11307
rect 16452 11248 17924 11307
rect 18280 11248 19752 11307
rect 20108 11248 21580 11307
rect 1630 11214 1708 11225
rect 3458 11214 3536 11225
rect 5286 11214 5364 11225
rect 7114 11214 7192 11225
rect 8942 11214 9020 11225
rect 10770 11214 10848 11225
rect 12598 11214 12676 11225
rect 14426 11214 14504 11225
rect 16254 11214 16332 11225
rect 18082 11214 18160 11225
rect 19910 11214 19988 11225
rect 21738 11214 21816 11225
rect 1488 11198 1708 11214
rect 1488 10822 1630 11198
rect 1488 10806 1708 10822
rect 3316 11198 3536 11214
rect 3316 10822 3458 11198
rect 3316 10806 3536 10822
rect 5144 11198 5364 11214
rect 5144 10822 5286 11198
rect 5144 10806 5364 10822
rect 6972 11198 7192 11214
rect 6972 10822 7114 11198
rect 6972 10806 7192 10822
rect 8800 11198 9020 11214
rect 8800 10822 8942 11198
rect 8800 10806 9020 10822
rect 10628 11198 10848 11214
rect 10628 10822 10770 11198
rect 10628 10806 10848 10822
rect 12456 11198 12676 11214
rect 12456 10822 12598 11198
rect 12456 10806 12676 10822
rect 14284 11198 14504 11214
rect 14284 10822 14426 11198
rect 14284 10806 14504 10822
rect 16112 11198 16332 11214
rect 16112 10822 16254 11198
rect 16112 10806 16332 10822
rect 17940 11198 18160 11214
rect 17940 10822 18082 11198
rect 17940 10806 18160 10822
rect 19768 11198 19988 11214
rect 19768 10822 19910 11198
rect 19768 10806 19988 10822
rect 21596 11198 21816 11214
rect 21596 10822 21738 11198
rect 21596 10806 21816 10822
rect 1630 10795 1708 10806
rect 3458 10795 3536 10806
rect 5286 10795 5364 10806
rect 7114 10795 7192 10806
rect 8942 10795 9020 10806
rect 10770 10795 10848 10806
rect 12598 10795 12676 10806
rect 14426 10795 14504 10806
rect 16254 10795 16332 10806
rect 18082 10795 18160 10806
rect 19910 10795 19988 10806
rect 21738 10795 21816 10806
rect 0 10713 1490 10772
rect 1828 10713 3318 10772
rect 3656 10713 5146 10772
rect 5484 10713 6974 10772
rect 7312 10713 8802 10772
rect 9140 10713 10630 10772
rect 10968 10713 12458 10772
rect 12796 10713 14286 10772
rect 14624 10713 16114 10772
rect 16452 10713 17942 10772
rect 18280 10713 19770 10772
rect 20108 10713 21598 10772
rect 0 10534 1472 10593
rect 1828 10534 3300 10593
rect 3656 10534 5128 10593
rect 5484 10534 6956 10593
rect 7312 10534 8784 10593
rect 9140 10534 10612 10593
rect 10968 10534 12440 10593
rect 12796 10534 14268 10593
rect 14624 10534 16096 10593
rect 16452 10534 17924 10593
rect 18280 10534 19752 10593
rect 20108 10534 21580 10593
rect 1630 10500 1708 10511
rect 3458 10500 3536 10511
rect 5286 10500 5364 10511
rect 7114 10500 7192 10511
rect 8942 10500 9020 10511
rect 10770 10500 10848 10511
rect 12598 10500 12676 10511
rect 14426 10500 14504 10511
rect 16254 10500 16332 10511
rect 18082 10500 18160 10511
rect 19910 10500 19988 10511
rect 21738 10500 21816 10511
rect 1488 10484 1708 10500
rect 1488 10108 1630 10484
rect 1488 10092 1708 10108
rect 3316 10484 3536 10500
rect 3316 10108 3458 10484
rect 3316 10092 3536 10108
rect 5144 10484 5364 10500
rect 5144 10108 5286 10484
rect 5144 10092 5364 10108
rect 6972 10484 7192 10500
rect 6972 10108 7114 10484
rect 6972 10092 7192 10108
rect 8800 10484 9020 10500
rect 8800 10108 8942 10484
rect 8800 10092 9020 10108
rect 10628 10484 10848 10500
rect 10628 10108 10770 10484
rect 10628 10092 10848 10108
rect 12456 10484 12676 10500
rect 12456 10108 12598 10484
rect 12456 10092 12676 10108
rect 14284 10484 14504 10500
rect 14284 10108 14426 10484
rect 14284 10092 14504 10108
rect 16112 10484 16332 10500
rect 16112 10108 16254 10484
rect 16112 10092 16332 10108
rect 17940 10484 18160 10500
rect 17940 10108 18082 10484
rect 17940 10092 18160 10108
rect 19768 10484 19988 10500
rect 19768 10108 19910 10484
rect 19768 10092 19988 10108
rect 21596 10484 21816 10500
rect 21596 10108 21738 10484
rect 21596 10092 21816 10108
rect 1630 10081 1708 10092
rect 3458 10081 3536 10092
rect 5286 10081 5364 10092
rect 7114 10081 7192 10092
rect 8942 10081 9020 10092
rect 10770 10081 10848 10092
rect 12598 10081 12676 10092
rect 14426 10081 14504 10092
rect 16254 10081 16332 10092
rect 18082 10081 18160 10092
rect 19910 10081 19988 10092
rect 21738 10081 21816 10092
rect 0 9999 1490 10058
rect 1828 9999 3318 10058
rect 3656 9999 5146 10058
rect 5484 9999 6974 10058
rect 7312 9999 8802 10058
rect 9140 9999 10630 10058
rect 10968 9999 12458 10058
rect 12796 9999 14286 10058
rect 14624 9999 16114 10058
rect 16452 9999 17942 10058
rect 18280 9999 19770 10058
rect 20108 9999 21598 10058
rect 0 9820 1472 9879
rect 1828 9820 3300 9879
rect 3656 9820 5128 9879
rect 5484 9820 6956 9879
rect 7312 9820 8784 9879
rect 9140 9820 10612 9879
rect 10968 9820 12440 9879
rect 12796 9820 14268 9879
rect 14624 9820 16096 9879
rect 16452 9820 17924 9879
rect 18280 9820 19752 9879
rect 20108 9820 21580 9879
rect 1630 9786 1708 9797
rect 3458 9786 3536 9797
rect 5286 9786 5364 9797
rect 7114 9786 7192 9797
rect 8942 9786 9020 9797
rect 10770 9786 10848 9797
rect 12598 9786 12676 9797
rect 14426 9786 14504 9797
rect 16254 9786 16332 9797
rect 18082 9786 18160 9797
rect 19910 9786 19988 9797
rect 21738 9786 21816 9797
rect 1488 9770 1708 9786
rect 1488 9394 1630 9770
rect 1488 9378 1708 9394
rect 3316 9770 3536 9786
rect 3316 9394 3458 9770
rect 3316 9378 3536 9394
rect 5144 9770 5364 9786
rect 5144 9394 5286 9770
rect 5144 9378 5364 9394
rect 6972 9770 7192 9786
rect 6972 9394 7114 9770
rect 6972 9378 7192 9394
rect 8800 9770 9020 9786
rect 8800 9394 8942 9770
rect 8800 9378 9020 9394
rect 10628 9770 10848 9786
rect 10628 9394 10770 9770
rect 10628 9378 10848 9394
rect 12456 9770 12676 9786
rect 12456 9394 12598 9770
rect 12456 9378 12676 9394
rect 14284 9770 14504 9786
rect 14284 9394 14426 9770
rect 14284 9378 14504 9394
rect 16112 9770 16332 9786
rect 16112 9394 16254 9770
rect 16112 9378 16332 9394
rect 17940 9770 18160 9786
rect 17940 9394 18082 9770
rect 17940 9378 18160 9394
rect 19768 9770 19988 9786
rect 19768 9394 19910 9770
rect 19768 9378 19988 9394
rect 21596 9770 21816 9786
rect 21596 9394 21738 9770
rect 21596 9378 21816 9394
rect 1630 9367 1708 9378
rect 3458 9367 3536 9378
rect 5286 9367 5364 9378
rect 7114 9367 7192 9378
rect 8942 9367 9020 9378
rect 10770 9367 10848 9378
rect 12598 9367 12676 9378
rect 14426 9367 14504 9378
rect 16254 9367 16332 9378
rect 18082 9367 18160 9378
rect 19910 9367 19988 9378
rect 21738 9367 21816 9378
rect 0 9285 1490 9344
rect 1828 9285 3318 9344
rect 3656 9285 5146 9344
rect 5484 9285 6974 9344
rect 7312 9285 8802 9344
rect 9140 9285 10630 9344
rect 10968 9285 12458 9344
rect 12796 9285 14286 9344
rect 14624 9285 16114 9344
rect 16452 9285 17942 9344
rect 18280 9285 19770 9344
rect 20108 9285 21598 9344
rect 0 9106 1472 9165
rect 1828 9106 3300 9165
rect 3656 9106 5128 9165
rect 5484 9106 6956 9165
rect 7312 9106 8784 9165
rect 9140 9106 10612 9165
rect 10968 9106 12440 9165
rect 12796 9106 14268 9165
rect 14624 9106 16096 9165
rect 16452 9106 17924 9165
rect 18280 9106 19752 9165
rect 20108 9106 21580 9165
rect 1630 9072 1708 9083
rect 3458 9072 3536 9083
rect 5286 9072 5364 9083
rect 7114 9072 7192 9083
rect 8942 9072 9020 9083
rect 10770 9072 10848 9083
rect 12598 9072 12676 9083
rect 14426 9072 14504 9083
rect 16254 9072 16332 9083
rect 18082 9072 18160 9083
rect 19910 9072 19988 9083
rect 21738 9072 21816 9083
rect 1488 9056 1708 9072
rect 1488 8680 1630 9056
rect 1488 8664 1708 8680
rect 3316 9056 3536 9072
rect 3316 8680 3458 9056
rect 3316 8664 3536 8680
rect 5144 9056 5364 9072
rect 5144 8680 5286 9056
rect 5144 8664 5364 8680
rect 6972 9056 7192 9072
rect 6972 8680 7114 9056
rect 6972 8664 7192 8680
rect 8800 9056 9020 9072
rect 8800 8680 8942 9056
rect 8800 8664 9020 8680
rect 10628 9056 10848 9072
rect 10628 8680 10770 9056
rect 10628 8664 10848 8680
rect 12456 9056 12676 9072
rect 12456 8680 12598 9056
rect 12456 8664 12676 8680
rect 14284 9056 14504 9072
rect 14284 8680 14426 9056
rect 14284 8664 14504 8680
rect 16112 9056 16332 9072
rect 16112 8680 16254 9056
rect 16112 8664 16332 8680
rect 17940 9056 18160 9072
rect 17940 8680 18082 9056
rect 17940 8664 18160 8680
rect 19768 9056 19988 9072
rect 19768 8680 19910 9056
rect 19768 8664 19988 8680
rect 21596 9056 21816 9072
rect 21596 8680 21738 9056
rect 21596 8664 21816 8680
rect 1630 8653 1708 8664
rect 3458 8653 3536 8664
rect 5286 8653 5364 8664
rect 7114 8653 7192 8664
rect 8942 8653 9020 8664
rect 10770 8653 10848 8664
rect 12598 8653 12676 8664
rect 14426 8653 14504 8664
rect 16254 8653 16332 8664
rect 18082 8653 18160 8664
rect 19910 8653 19988 8664
rect 21738 8653 21816 8664
rect 0 8571 1490 8630
rect 1828 8571 3318 8630
rect 3656 8571 5146 8630
rect 5484 8571 6974 8630
rect 7312 8571 8802 8630
rect 9140 8571 10630 8630
rect 10968 8571 12458 8630
rect 12796 8571 14286 8630
rect 14624 8571 16114 8630
rect 16452 8571 17942 8630
rect 18280 8571 19770 8630
rect 20108 8571 21598 8630
rect 0 8392 1472 8451
rect 1828 8392 3300 8451
rect 3656 8392 5128 8451
rect 5484 8392 6956 8451
rect 7312 8392 8784 8451
rect 9140 8392 10612 8451
rect 10968 8392 12440 8451
rect 12796 8392 14268 8451
rect 14624 8392 16096 8451
rect 16452 8392 17924 8451
rect 18280 8392 19752 8451
rect 20108 8392 21580 8451
rect 1630 8358 1708 8369
rect 3458 8358 3536 8369
rect 5286 8358 5364 8369
rect 7114 8358 7192 8369
rect 8942 8358 9020 8369
rect 10770 8358 10848 8369
rect 12598 8358 12676 8369
rect 14426 8358 14504 8369
rect 16254 8358 16332 8369
rect 18082 8358 18160 8369
rect 19910 8358 19988 8369
rect 21738 8358 21816 8369
rect 1488 8342 1708 8358
rect 1488 7966 1630 8342
rect 1488 7950 1708 7966
rect 3316 8342 3536 8358
rect 3316 7966 3458 8342
rect 3316 7950 3536 7966
rect 5144 8342 5364 8358
rect 5144 7966 5286 8342
rect 5144 7950 5364 7966
rect 6972 8342 7192 8358
rect 6972 7966 7114 8342
rect 6972 7950 7192 7966
rect 8800 8342 9020 8358
rect 8800 7966 8942 8342
rect 8800 7950 9020 7966
rect 10628 8342 10848 8358
rect 10628 7966 10770 8342
rect 10628 7950 10848 7966
rect 12456 8342 12676 8358
rect 12456 7966 12598 8342
rect 12456 7950 12676 7966
rect 14284 8342 14504 8358
rect 14284 7966 14426 8342
rect 14284 7950 14504 7966
rect 16112 8342 16332 8358
rect 16112 7966 16254 8342
rect 16112 7950 16332 7966
rect 17940 8342 18160 8358
rect 17940 7966 18082 8342
rect 17940 7950 18160 7966
rect 19768 8342 19988 8358
rect 19768 7966 19910 8342
rect 19768 7950 19988 7966
rect 21596 8342 21816 8358
rect 21596 7966 21738 8342
rect 21596 7950 21816 7966
rect 1630 7939 1708 7950
rect 3458 7939 3536 7950
rect 5286 7939 5364 7950
rect 7114 7939 7192 7950
rect 8942 7939 9020 7950
rect 10770 7939 10848 7950
rect 12598 7939 12676 7950
rect 14426 7939 14504 7950
rect 16254 7939 16332 7950
rect 18082 7939 18160 7950
rect 19910 7939 19988 7950
rect 21738 7939 21816 7950
rect 0 7857 1490 7916
rect 1828 7857 3318 7916
rect 3656 7857 5146 7916
rect 5484 7857 6974 7916
rect 7312 7857 8802 7916
rect 9140 7857 10630 7916
rect 10968 7857 12458 7916
rect 12796 7857 14286 7916
rect 14624 7857 16114 7916
rect 16452 7857 17942 7916
rect 18280 7857 19770 7916
rect 20108 7857 21598 7916
rect 0 7678 1472 7737
rect 1828 7678 3300 7737
rect 3656 7678 5128 7737
rect 5484 7678 6956 7737
rect 7312 7678 8784 7737
rect 9140 7678 10612 7737
rect 10968 7678 12440 7737
rect 12796 7678 14268 7737
rect 14624 7678 16096 7737
rect 16452 7678 17924 7737
rect 18280 7678 19752 7737
rect 20108 7678 21580 7737
rect 1630 7644 1708 7655
rect 3458 7644 3536 7655
rect 5286 7644 5364 7655
rect 7114 7644 7192 7655
rect 8942 7644 9020 7655
rect 10770 7644 10848 7655
rect 12598 7644 12676 7655
rect 14426 7644 14504 7655
rect 16254 7644 16332 7655
rect 18082 7644 18160 7655
rect 19910 7644 19988 7655
rect 21738 7644 21816 7655
rect 1488 7628 1708 7644
rect 1488 7252 1630 7628
rect 1488 7236 1708 7252
rect 3316 7628 3536 7644
rect 3316 7252 3458 7628
rect 3316 7236 3536 7252
rect 5144 7628 5364 7644
rect 5144 7252 5286 7628
rect 5144 7236 5364 7252
rect 6972 7628 7192 7644
rect 6972 7252 7114 7628
rect 6972 7236 7192 7252
rect 8800 7628 9020 7644
rect 8800 7252 8942 7628
rect 8800 7236 9020 7252
rect 10628 7628 10848 7644
rect 10628 7252 10770 7628
rect 10628 7236 10848 7252
rect 12456 7628 12676 7644
rect 12456 7252 12598 7628
rect 12456 7236 12676 7252
rect 14284 7628 14504 7644
rect 14284 7252 14426 7628
rect 14284 7236 14504 7252
rect 16112 7628 16332 7644
rect 16112 7252 16254 7628
rect 16112 7236 16332 7252
rect 17940 7628 18160 7644
rect 17940 7252 18082 7628
rect 17940 7236 18160 7252
rect 19768 7628 19988 7644
rect 19768 7252 19910 7628
rect 19768 7236 19988 7252
rect 21596 7628 21816 7644
rect 21596 7252 21738 7628
rect 21596 7236 21816 7252
rect 1630 7225 1708 7236
rect 3458 7225 3536 7236
rect 5286 7225 5364 7236
rect 7114 7225 7192 7236
rect 8942 7225 9020 7236
rect 10770 7225 10848 7236
rect 12598 7225 12676 7236
rect 14426 7225 14504 7236
rect 16254 7225 16332 7236
rect 18082 7225 18160 7236
rect 19910 7225 19988 7236
rect 21738 7225 21816 7236
rect 0 7143 1490 7202
rect 1828 7143 3318 7202
rect 3656 7143 5146 7202
rect 5484 7143 6974 7202
rect 7312 7143 8802 7202
rect 9140 7143 10630 7202
rect 10968 7143 12458 7202
rect 12796 7143 14286 7202
rect 14624 7143 16114 7202
rect 16452 7143 17942 7202
rect 18280 7143 19770 7202
rect 20108 7143 21598 7202
rect 0 6964 1472 7023
rect 1828 6964 3300 7023
rect 3656 6964 5128 7023
rect 5484 6964 6956 7023
rect 7312 6964 8784 7023
rect 9140 6964 10612 7023
rect 10968 6964 12440 7023
rect 12796 6964 14268 7023
rect 14624 6964 16096 7023
rect 16452 6964 17924 7023
rect 18280 6964 19752 7023
rect 20108 6964 21580 7023
rect 1630 6930 1708 6941
rect 3458 6930 3536 6941
rect 5286 6930 5364 6941
rect 7114 6930 7192 6941
rect 8942 6930 9020 6941
rect 10770 6930 10848 6941
rect 12598 6930 12676 6941
rect 14426 6930 14504 6941
rect 16254 6930 16332 6941
rect 18082 6930 18160 6941
rect 19910 6930 19988 6941
rect 21738 6930 21816 6941
rect 1488 6914 1708 6930
rect 1488 6538 1630 6914
rect 1488 6522 1708 6538
rect 3316 6914 3536 6930
rect 3316 6538 3458 6914
rect 3316 6522 3536 6538
rect 5144 6914 5364 6930
rect 5144 6538 5286 6914
rect 5144 6522 5364 6538
rect 6972 6914 7192 6930
rect 6972 6538 7114 6914
rect 6972 6522 7192 6538
rect 8800 6914 9020 6930
rect 8800 6538 8942 6914
rect 8800 6522 9020 6538
rect 10628 6914 10848 6930
rect 10628 6538 10770 6914
rect 10628 6522 10848 6538
rect 12456 6914 12676 6930
rect 12456 6538 12598 6914
rect 12456 6522 12676 6538
rect 14284 6914 14504 6930
rect 14284 6538 14426 6914
rect 14284 6522 14504 6538
rect 16112 6914 16332 6930
rect 16112 6538 16254 6914
rect 16112 6522 16332 6538
rect 17940 6914 18160 6930
rect 17940 6538 18082 6914
rect 17940 6522 18160 6538
rect 19768 6914 19988 6930
rect 19768 6538 19910 6914
rect 19768 6522 19988 6538
rect 21596 6914 21816 6930
rect 21596 6538 21738 6914
rect 21596 6522 21816 6538
rect 1630 6511 1708 6522
rect 3458 6511 3536 6522
rect 5286 6511 5364 6522
rect 7114 6511 7192 6522
rect 8942 6511 9020 6522
rect 10770 6511 10848 6522
rect 12598 6511 12676 6522
rect 14426 6511 14504 6522
rect 16254 6511 16332 6522
rect 18082 6511 18160 6522
rect 19910 6511 19988 6522
rect 21738 6511 21816 6522
rect 0 6429 1490 6488
rect 1828 6429 3318 6488
rect 3656 6429 5146 6488
rect 5484 6429 6974 6488
rect 7312 6429 8802 6488
rect 9140 6429 10630 6488
rect 10968 6429 12458 6488
rect 12796 6429 14286 6488
rect 14624 6429 16114 6488
rect 16452 6429 17942 6488
rect 18280 6429 19770 6488
rect 20108 6429 21598 6488
rect 0 6250 1472 6309
rect 1828 6250 3300 6309
rect 3656 6250 5128 6309
rect 5484 6250 6956 6309
rect 7312 6250 8784 6309
rect 9140 6250 10612 6309
rect 10968 6250 12440 6309
rect 12796 6250 14268 6309
rect 14624 6250 16096 6309
rect 16452 6250 17924 6309
rect 18280 6250 19752 6309
rect 20108 6250 21580 6309
rect 1630 6216 1708 6227
rect 3458 6216 3536 6227
rect 5286 6216 5364 6227
rect 7114 6216 7192 6227
rect 8942 6216 9020 6227
rect 10770 6216 10848 6227
rect 12598 6216 12676 6227
rect 14426 6216 14504 6227
rect 16254 6216 16332 6227
rect 18082 6216 18160 6227
rect 19910 6216 19988 6227
rect 21738 6216 21816 6227
rect 1488 6200 1708 6216
rect 1488 5824 1630 6200
rect 1488 5808 1708 5824
rect 3316 6200 3536 6216
rect 3316 5824 3458 6200
rect 3316 5808 3536 5824
rect 5144 6200 5364 6216
rect 5144 5824 5286 6200
rect 5144 5808 5364 5824
rect 6972 6200 7192 6216
rect 6972 5824 7114 6200
rect 6972 5808 7192 5824
rect 8800 6200 9020 6216
rect 8800 5824 8942 6200
rect 8800 5808 9020 5824
rect 10628 6200 10848 6216
rect 10628 5824 10770 6200
rect 10628 5808 10848 5824
rect 12456 6200 12676 6216
rect 12456 5824 12598 6200
rect 12456 5808 12676 5824
rect 14284 6200 14504 6216
rect 14284 5824 14426 6200
rect 14284 5808 14504 5824
rect 16112 6200 16332 6216
rect 16112 5824 16254 6200
rect 16112 5808 16332 5824
rect 17940 6200 18160 6216
rect 17940 5824 18082 6200
rect 17940 5808 18160 5824
rect 19768 6200 19988 6216
rect 19768 5824 19910 6200
rect 19768 5808 19988 5824
rect 21596 6200 21816 6216
rect 21596 5824 21738 6200
rect 21596 5808 21816 5824
rect 1630 5797 1708 5808
rect 3458 5797 3536 5808
rect 5286 5797 5364 5808
rect 7114 5797 7192 5808
rect 8942 5797 9020 5808
rect 10770 5797 10848 5808
rect 12598 5797 12676 5808
rect 14426 5797 14504 5808
rect 16254 5797 16332 5808
rect 18082 5797 18160 5808
rect 19910 5797 19988 5808
rect 21738 5797 21816 5808
rect 0 5715 1490 5774
rect 1828 5715 3318 5774
rect 3656 5715 5146 5774
rect 5484 5715 6974 5774
rect 7312 5715 8802 5774
rect 9140 5715 10630 5774
rect 10968 5715 12458 5774
rect 12796 5715 14286 5774
rect 14624 5715 16114 5774
rect 16452 5715 17942 5774
rect 18280 5715 19770 5774
rect 20108 5715 21598 5774
rect 0 5536 1472 5595
rect 1828 5536 3300 5595
rect 3656 5536 5128 5595
rect 5484 5536 6956 5595
rect 7312 5536 8784 5595
rect 9140 5536 10612 5595
rect 10968 5536 12440 5595
rect 12796 5536 14268 5595
rect 14624 5536 16096 5595
rect 16452 5536 17924 5595
rect 18280 5536 19752 5595
rect 20108 5536 21580 5595
rect 1630 5502 1708 5513
rect 3458 5502 3536 5513
rect 5286 5502 5364 5513
rect 7114 5502 7192 5513
rect 8942 5502 9020 5513
rect 10770 5502 10848 5513
rect 12598 5502 12676 5513
rect 14426 5502 14504 5513
rect 16254 5502 16332 5513
rect 18082 5502 18160 5513
rect 19910 5502 19988 5513
rect 21738 5502 21816 5513
rect 1488 5486 1708 5502
rect 1488 5110 1630 5486
rect 1488 5094 1708 5110
rect 3316 5486 3536 5502
rect 3316 5110 3458 5486
rect 3316 5094 3536 5110
rect 5144 5486 5364 5502
rect 5144 5110 5286 5486
rect 5144 5094 5364 5110
rect 6972 5486 7192 5502
rect 6972 5110 7114 5486
rect 6972 5094 7192 5110
rect 8800 5486 9020 5502
rect 8800 5110 8942 5486
rect 8800 5094 9020 5110
rect 10628 5486 10848 5502
rect 10628 5110 10770 5486
rect 10628 5094 10848 5110
rect 12456 5486 12676 5502
rect 12456 5110 12598 5486
rect 12456 5094 12676 5110
rect 14284 5486 14504 5502
rect 14284 5110 14426 5486
rect 14284 5094 14504 5110
rect 16112 5486 16332 5502
rect 16112 5110 16254 5486
rect 16112 5094 16332 5110
rect 17940 5486 18160 5502
rect 17940 5110 18082 5486
rect 17940 5094 18160 5110
rect 19768 5486 19988 5502
rect 19768 5110 19910 5486
rect 19768 5094 19988 5110
rect 21596 5486 21816 5502
rect 21596 5110 21738 5486
rect 21596 5094 21816 5110
rect 1630 5083 1708 5094
rect 3458 5083 3536 5094
rect 5286 5083 5364 5094
rect 7114 5083 7192 5094
rect 8942 5083 9020 5094
rect 10770 5083 10848 5094
rect 12598 5083 12676 5094
rect 14426 5083 14504 5094
rect 16254 5083 16332 5094
rect 18082 5083 18160 5094
rect 19910 5083 19988 5094
rect 21738 5083 21816 5094
rect 0 5001 1490 5060
rect 1828 5001 3318 5060
rect 3656 5001 5146 5060
rect 5484 5001 6974 5060
rect 7312 5001 8802 5060
rect 9140 5001 10630 5060
rect 10968 5001 12458 5060
rect 12796 5001 14286 5060
rect 14624 5001 16114 5060
rect 16452 5001 17942 5060
rect 18280 5001 19770 5060
rect 20108 5001 21598 5060
rect 0 4822 1472 4881
rect 1828 4822 3300 4881
rect 3656 4822 5128 4881
rect 5484 4822 6956 4881
rect 7312 4822 8784 4881
rect 9140 4822 10612 4881
rect 10968 4822 12440 4881
rect 12796 4822 14268 4881
rect 14624 4822 16096 4881
rect 16452 4822 17924 4881
rect 18280 4822 19752 4881
rect 20108 4822 21580 4881
rect 1630 4788 1708 4799
rect 3458 4788 3536 4799
rect 5286 4788 5364 4799
rect 7114 4788 7192 4799
rect 8942 4788 9020 4799
rect 10770 4788 10848 4799
rect 12598 4788 12676 4799
rect 14426 4788 14504 4799
rect 16254 4788 16332 4799
rect 18082 4788 18160 4799
rect 19910 4788 19988 4799
rect 21738 4788 21816 4799
rect 1488 4772 1708 4788
rect 1488 4396 1630 4772
rect 1488 4380 1708 4396
rect 3316 4772 3536 4788
rect 3316 4396 3458 4772
rect 3316 4380 3536 4396
rect 5144 4772 5364 4788
rect 5144 4396 5286 4772
rect 5144 4380 5364 4396
rect 6972 4772 7192 4788
rect 6972 4396 7114 4772
rect 6972 4380 7192 4396
rect 8800 4772 9020 4788
rect 8800 4396 8942 4772
rect 8800 4380 9020 4396
rect 10628 4772 10848 4788
rect 10628 4396 10770 4772
rect 10628 4380 10848 4396
rect 12456 4772 12676 4788
rect 12456 4396 12598 4772
rect 12456 4380 12676 4396
rect 14284 4772 14504 4788
rect 14284 4396 14426 4772
rect 14284 4380 14504 4396
rect 16112 4772 16332 4788
rect 16112 4396 16254 4772
rect 16112 4380 16332 4396
rect 17940 4772 18160 4788
rect 17940 4396 18082 4772
rect 17940 4380 18160 4396
rect 19768 4772 19988 4788
rect 19768 4396 19910 4772
rect 19768 4380 19988 4396
rect 21596 4772 21816 4788
rect 21596 4396 21738 4772
rect 21596 4380 21816 4396
rect 1630 4369 1708 4380
rect 3458 4369 3536 4380
rect 5286 4369 5364 4380
rect 7114 4369 7192 4380
rect 8942 4369 9020 4380
rect 10770 4369 10848 4380
rect 12598 4369 12676 4380
rect 14426 4369 14504 4380
rect 16254 4369 16332 4380
rect 18082 4369 18160 4380
rect 19910 4369 19988 4380
rect 21738 4369 21816 4380
rect 0 4287 1490 4346
rect 1828 4287 3318 4346
rect 3656 4287 5146 4346
rect 5484 4287 6974 4346
rect 7312 4287 8802 4346
rect 9140 4287 10630 4346
rect 10968 4287 12458 4346
rect 12796 4287 14286 4346
rect 14624 4287 16114 4346
rect 16452 4287 17942 4346
rect 18280 4287 19770 4346
rect 20108 4287 21598 4346
rect 0 4108 1472 4167
rect 1828 4108 3300 4167
rect 3656 4108 5128 4167
rect 5484 4108 6956 4167
rect 7312 4108 8784 4167
rect 9140 4108 10612 4167
rect 10968 4108 12440 4167
rect 12796 4108 14268 4167
rect 14624 4108 16096 4167
rect 16452 4108 17924 4167
rect 18280 4108 19752 4167
rect 20108 4108 21580 4167
rect 1630 4074 1708 4085
rect 3458 4074 3536 4085
rect 5286 4074 5364 4085
rect 7114 4074 7192 4085
rect 8942 4074 9020 4085
rect 10770 4074 10848 4085
rect 12598 4074 12676 4085
rect 14426 4074 14504 4085
rect 16254 4074 16332 4085
rect 18082 4074 18160 4085
rect 19910 4074 19988 4085
rect 21738 4074 21816 4085
rect 1488 4058 1708 4074
rect 1488 3682 1630 4058
rect 1488 3666 1708 3682
rect 3316 4058 3536 4074
rect 3316 3682 3458 4058
rect 3316 3666 3536 3682
rect 5144 4058 5364 4074
rect 5144 3682 5286 4058
rect 5144 3666 5364 3682
rect 6972 4058 7192 4074
rect 6972 3682 7114 4058
rect 6972 3666 7192 3682
rect 8800 4058 9020 4074
rect 8800 3682 8942 4058
rect 8800 3666 9020 3682
rect 10628 4058 10848 4074
rect 10628 3682 10770 4058
rect 10628 3666 10848 3682
rect 12456 4058 12676 4074
rect 12456 3682 12598 4058
rect 12456 3666 12676 3682
rect 14284 4058 14504 4074
rect 14284 3682 14426 4058
rect 14284 3666 14504 3682
rect 16112 4058 16332 4074
rect 16112 3682 16254 4058
rect 16112 3666 16332 3682
rect 17940 4058 18160 4074
rect 17940 3682 18082 4058
rect 17940 3666 18160 3682
rect 19768 4058 19988 4074
rect 19768 3682 19910 4058
rect 19768 3666 19988 3682
rect 21596 4058 21816 4074
rect 21596 3682 21738 4058
rect 21596 3666 21816 3682
rect 1630 3655 1708 3666
rect 3458 3655 3536 3666
rect 5286 3655 5364 3666
rect 7114 3655 7192 3666
rect 8942 3655 9020 3666
rect 10770 3655 10848 3666
rect 12598 3655 12676 3666
rect 14426 3655 14504 3666
rect 16254 3655 16332 3666
rect 18082 3655 18160 3666
rect 19910 3655 19988 3666
rect 21738 3655 21816 3666
rect 0 3573 1490 3632
rect 1828 3573 3318 3632
rect 3656 3573 5146 3632
rect 5484 3573 6974 3632
rect 7312 3573 8802 3632
rect 9140 3573 10630 3632
rect 10968 3573 12458 3632
rect 12796 3573 14286 3632
rect 14624 3573 16114 3632
rect 16452 3573 17942 3632
rect 18280 3573 19770 3632
rect 20108 3573 21598 3632
rect 0 3394 1472 3453
rect 1828 3394 3300 3453
rect 3656 3394 5128 3453
rect 5484 3394 6956 3453
rect 7312 3394 8784 3453
rect 9140 3394 10612 3453
rect 10968 3394 12440 3453
rect 12796 3394 14268 3453
rect 14624 3394 16096 3453
rect 16452 3394 17924 3453
rect 18280 3394 19752 3453
rect 20108 3394 21580 3453
rect 1630 3360 1708 3371
rect 3458 3360 3536 3371
rect 5286 3360 5364 3371
rect 7114 3360 7192 3371
rect 8942 3360 9020 3371
rect 10770 3360 10848 3371
rect 12598 3360 12676 3371
rect 14426 3360 14504 3371
rect 16254 3360 16332 3371
rect 18082 3360 18160 3371
rect 19910 3360 19988 3371
rect 21738 3360 21816 3371
rect 1488 3344 1708 3360
rect 1488 2968 1630 3344
rect 1488 2952 1708 2968
rect 3316 3344 3536 3360
rect 3316 2968 3458 3344
rect 3316 2952 3536 2968
rect 5144 3344 5364 3360
rect 5144 2968 5286 3344
rect 5144 2952 5364 2968
rect 6972 3344 7192 3360
rect 6972 2968 7114 3344
rect 6972 2952 7192 2968
rect 8800 3344 9020 3360
rect 8800 2968 8942 3344
rect 8800 2952 9020 2968
rect 10628 3344 10848 3360
rect 10628 2968 10770 3344
rect 10628 2952 10848 2968
rect 12456 3344 12676 3360
rect 12456 2968 12598 3344
rect 12456 2952 12676 2968
rect 14284 3344 14504 3360
rect 14284 2968 14426 3344
rect 14284 2952 14504 2968
rect 16112 3344 16332 3360
rect 16112 2968 16254 3344
rect 16112 2952 16332 2968
rect 17940 3344 18160 3360
rect 17940 2968 18082 3344
rect 17940 2952 18160 2968
rect 19768 3344 19988 3360
rect 19768 2968 19910 3344
rect 19768 2952 19988 2968
rect 21596 3344 21816 3360
rect 21596 2968 21738 3344
rect 21596 2952 21816 2968
rect 1630 2941 1708 2952
rect 3458 2941 3536 2952
rect 5286 2941 5364 2952
rect 7114 2941 7192 2952
rect 8942 2941 9020 2952
rect 10770 2941 10848 2952
rect 12598 2941 12676 2952
rect 14426 2941 14504 2952
rect 16254 2941 16332 2952
rect 18082 2941 18160 2952
rect 19910 2941 19988 2952
rect 21738 2941 21816 2952
rect 0 2859 1490 2918
rect 1828 2859 3318 2918
rect 3656 2859 5146 2918
rect 5484 2859 6974 2918
rect 7312 2859 8802 2918
rect 9140 2859 10630 2918
rect 10968 2859 12458 2918
rect 12796 2859 14286 2918
rect 14624 2859 16114 2918
rect 16452 2859 17942 2918
rect 18280 2859 19770 2918
rect 20108 2859 21598 2918
rect 0 2680 1472 2739
rect 1828 2680 3300 2739
rect 3656 2680 5128 2739
rect 5484 2680 6956 2739
rect 7312 2680 8784 2739
rect 9140 2680 10612 2739
rect 10968 2680 12440 2739
rect 12796 2680 14268 2739
rect 14624 2680 16096 2739
rect 16452 2680 17924 2739
rect 18280 2680 19752 2739
rect 20108 2680 21580 2739
rect 1630 2646 1708 2657
rect 3458 2646 3536 2657
rect 5286 2646 5364 2657
rect 7114 2646 7192 2657
rect 8942 2646 9020 2657
rect 10770 2646 10848 2657
rect 12598 2646 12676 2657
rect 14426 2646 14504 2657
rect 16254 2646 16332 2657
rect 18082 2646 18160 2657
rect 19910 2646 19988 2657
rect 21738 2646 21816 2657
rect 1488 2630 1708 2646
rect 1488 2254 1630 2630
rect 1488 2238 1708 2254
rect 3316 2630 3536 2646
rect 3316 2254 3458 2630
rect 3316 2238 3536 2254
rect 5144 2630 5364 2646
rect 5144 2254 5286 2630
rect 5144 2238 5364 2254
rect 6972 2630 7192 2646
rect 6972 2254 7114 2630
rect 6972 2238 7192 2254
rect 8800 2630 9020 2646
rect 8800 2254 8942 2630
rect 8800 2238 9020 2254
rect 10628 2630 10848 2646
rect 10628 2254 10770 2630
rect 10628 2238 10848 2254
rect 12456 2630 12676 2646
rect 12456 2254 12598 2630
rect 12456 2238 12676 2254
rect 14284 2630 14504 2646
rect 14284 2254 14426 2630
rect 14284 2238 14504 2254
rect 16112 2630 16332 2646
rect 16112 2254 16254 2630
rect 16112 2238 16332 2254
rect 17940 2630 18160 2646
rect 17940 2254 18082 2630
rect 17940 2238 18160 2254
rect 19768 2630 19988 2646
rect 19768 2254 19910 2630
rect 19768 2238 19988 2254
rect 21596 2630 21816 2646
rect 21596 2254 21738 2630
rect 21596 2238 21816 2254
rect 1630 2227 1708 2238
rect 3458 2227 3536 2238
rect 5286 2227 5364 2238
rect 7114 2227 7192 2238
rect 8942 2227 9020 2238
rect 10770 2227 10848 2238
rect 12598 2227 12676 2238
rect 14426 2227 14504 2238
rect 16254 2227 16332 2238
rect 18082 2227 18160 2238
rect 19910 2227 19988 2238
rect 21738 2227 21816 2238
rect 0 2145 1490 2204
rect 1828 2145 3318 2204
rect 3656 2145 5146 2204
rect 5484 2145 6974 2204
rect 7312 2145 8802 2204
rect 9140 2145 10630 2204
rect 10968 2145 12458 2204
rect 12796 2145 14286 2204
rect 14624 2145 16114 2204
rect 16452 2145 17942 2204
rect 18280 2145 19770 2204
rect 20108 2145 21598 2204
rect 0 1966 1472 2025
rect 1828 1966 3300 2025
rect 3656 1966 5128 2025
rect 5484 1966 6956 2025
rect 7312 1966 8784 2025
rect 9140 1966 10612 2025
rect 10968 1966 12440 2025
rect 12796 1966 14268 2025
rect 14624 1966 16096 2025
rect 16452 1966 17924 2025
rect 18280 1966 19752 2025
rect 20108 1966 21580 2025
rect 1630 1932 1708 1943
rect 3458 1932 3536 1943
rect 5286 1932 5364 1943
rect 7114 1932 7192 1943
rect 8942 1932 9020 1943
rect 10770 1932 10848 1943
rect 12598 1932 12676 1943
rect 14426 1932 14504 1943
rect 16254 1932 16332 1943
rect 18082 1932 18160 1943
rect 19910 1932 19988 1943
rect 21738 1932 21816 1943
rect 1488 1916 1708 1932
rect 1488 1540 1630 1916
rect 1488 1524 1708 1540
rect 3316 1916 3536 1932
rect 3316 1540 3458 1916
rect 3316 1524 3536 1540
rect 5144 1916 5364 1932
rect 5144 1540 5286 1916
rect 5144 1524 5364 1540
rect 6972 1916 7192 1932
rect 6972 1540 7114 1916
rect 6972 1524 7192 1540
rect 8800 1916 9020 1932
rect 8800 1540 8942 1916
rect 8800 1524 9020 1540
rect 10628 1916 10848 1932
rect 10628 1540 10770 1916
rect 10628 1524 10848 1540
rect 12456 1916 12676 1932
rect 12456 1540 12598 1916
rect 12456 1524 12676 1540
rect 14284 1916 14504 1932
rect 14284 1540 14426 1916
rect 14284 1524 14504 1540
rect 16112 1916 16332 1932
rect 16112 1540 16254 1916
rect 16112 1524 16332 1540
rect 17940 1916 18160 1932
rect 17940 1540 18082 1916
rect 17940 1524 18160 1540
rect 19768 1916 19988 1932
rect 19768 1540 19910 1916
rect 19768 1524 19988 1540
rect 21596 1916 21816 1932
rect 21596 1540 21738 1916
rect 21596 1524 21816 1540
rect 1630 1513 1708 1524
rect 3458 1513 3536 1524
rect 5286 1513 5364 1524
rect 7114 1513 7192 1524
rect 8942 1513 9020 1524
rect 10770 1513 10848 1524
rect 12598 1513 12676 1524
rect 14426 1513 14504 1524
rect 16254 1513 16332 1524
rect 18082 1513 18160 1524
rect 19910 1513 19988 1524
rect 21738 1513 21816 1524
rect 0 1431 1490 1490
rect 1828 1431 3318 1490
rect 3656 1431 5146 1490
rect 5484 1431 6974 1490
rect 7312 1431 8802 1490
rect 9140 1431 10630 1490
rect 10968 1431 12458 1490
rect 12796 1431 14286 1490
rect 14624 1431 16114 1490
rect 16452 1431 17942 1490
rect 18280 1431 19770 1490
rect 20108 1431 21598 1490
rect 0 1252 1472 1311
rect 1828 1252 3300 1311
rect 3656 1252 5128 1311
rect 5484 1252 6956 1311
rect 7312 1252 8784 1311
rect 9140 1252 10612 1311
rect 10968 1252 12440 1311
rect 12796 1252 14268 1311
rect 14624 1252 16096 1311
rect 16452 1252 17924 1311
rect 18280 1252 19752 1311
rect 20108 1252 21580 1311
rect 1630 1218 1708 1229
rect 3458 1218 3536 1229
rect 5286 1218 5364 1229
rect 7114 1218 7192 1229
rect 8942 1218 9020 1229
rect 10770 1218 10848 1229
rect 12598 1218 12676 1229
rect 14426 1218 14504 1229
rect 16254 1218 16332 1229
rect 18082 1218 18160 1229
rect 19910 1218 19988 1229
rect 21738 1218 21816 1229
rect 1488 1202 1708 1218
rect 1488 826 1630 1202
rect 1488 810 1708 826
rect 3316 1202 3536 1218
rect 3316 826 3458 1202
rect 3316 810 3536 826
rect 5144 1202 5364 1218
rect 5144 826 5286 1202
rect 5144 810 5364 826
rect 6972 1202 7192 1218
rect 6972 826 7114 1202
rect 6972 810 7192 826
rect 8800 1202 9020 1218
rect 8800 826 8942 1202
rect 8800 810 9020 826
rect 10628 1202 10848 1218
rect 10628 826 10770 1202
rect 10628 810 10848 826
rect 12456 1202 12676 1218
rect 12456 826 12598 1202
rect 12456 810 12676 826
rect 14284 1202 14504 1218
rect 14284 826 14426 1202
rect 14284 810 14504 826
rect 16112 1202 16332 1218
rect 16112 826 16254 1202
rect 16112 810 16332 826
rect 17940 1202 18160 1218
rect 17940 826 18082 1202
rect 17940 810 18160 826
rect 19768 1202 19988 1218
rect 19768 826 19910 1202
rect 19768 810 19988 826
rect 21596 1202 21816 1218
rect 21596 826 21738 1202
rect 21596 810 21816 826
rect 1630 799 1708 810
rect 3458 799 3536 810
rect 5286 799 5364 810
rect 7114 799 7192 810
rect 8942 799 9020 810
rect 10770 799 10848 810
rect 12598 799 12676 810
rect 14426 799 14504 810
rect 16254 799 16332 810
rect 18082 799 18160 810
rect 19910 799 19988 810
rect 21738 799 21816 810
rect 0 717 1490 776
rect 1828 717 3318 776
rect 3656 717 5146 776
rect 5484 717 6974 776
rect 7312 717 8802 776
rect 9140 717 10630 776
rect 10968 717 12458 776
rect 12796 717 14286 776
rect 14624 717 16114 776
rect 16452 717 17942 776
rect 18280 717 19770 776
rect 20108 717 21598 776
rect 0 538 1472 597
rect 1828 538 3300 597
rect 3656 538 5128 597
rect 5484 538 6956 597
rect 7312 538 8784 597
rect 9140 538 10612 597
rect 10968 538 12440 597
rect 12796 538 14268 597
rect 14624 538 16096 597
rect 16452 538 17924 597
rect 18280 538 19752 597
rect 20108 538 21580 597
rect 1630 504 1708 515
rect 3458 504 3536 515
rect 5286 504 5364 515
rect 7114 504 7192 515
rect 8942 504 9020 515
rect 10770 504 10848 515
rect 12598 504 12676 515
rect 14426 504 14504 515
rect 16254 504 16332 515
rect 18082 504 18160 515
rect 19910 504 19988 515
rect 21738 504 21816 515
rect 1488 488 1708 504
rect 1488 112 1630 488
rect 1488 96 1708 112
rect 3316 488 3536 504
rect 3316 112 3458 488
rect 3316 96 3536 112
rect 5144 488 5364 504
rect 5144 112 5286 488
rect 5144 96 5364 112
rect 6972 488 7192 504
rect 6972 112 7114 488
rect 6972 96 7192 112
rect 8800 488 9020 504
rect 8800 112 8942 488
rect 8800 96 9020 112
rect 10628 488 10848 504
rect 10628 112 10770 488
rect 10628 96 10848 112
rect 12456 488 12676 504
rect 12456 112 12598 488
rect 12456 96 12676 112
rect 14284 488 14504 504
rect 14284 112 14426 488
rect 14284 96 14504 112
rect 16112 488 16332 504
rect 16112 112 16254 488
rect 16112 96 16332 112
rect 17940 488 18160 504
rect 17940 112 18082 488
rect 17940 96 18160 112
rect 19768 488 19988 504
rect 19768 112 19910 488
rect 19768 96 19988 112
rect 21596 488 21816 504
rect 21596 112 21738 488
rect 21596 96 21816 112
rect 1630 85 1708 96
rect 3458 85 3536 96
rect 5286 85 5364 96
rect 7114 85 7192 96
rect 8942 85 9020 96
rect 10770 85 10848 96
rect 12598 85 12676 96
rect 14426 85 14504 96
rect 16254 85 16332 96
rect 18082 85 18160 96
rect 19910 85 19988 96
rect 21738 85 21816 96
rect 0 3 1490 62
rect 1828 3 3318 62
rect 3656 3 5146 62
rect 5484 3 6974 62
rect 7312 3 8802 62
rect 9140 3 10630 62
rect 10968 3 12458 62
rect 12796 3 14286 62
rect 14624 3 16114 62
rect 16452 3 17942 62
rect 18280 3 19770 62
rect 20108 3 21598 62
<< metal1 >>
rect 0 21244 1490 21303
rect 1828 21244 3318 21303
rect 3656 21244 5146 21303
rect 5484 21244 6974 21303
rect 7312 21244 8802 21303
rect 9140 21244 10630 21303
rect 10968 21244 12458 21303
rect 12796 21244 14286 21303
rect 14624 21244 16114 21303
rect 16452 21244 17942 21303
rect 18280 21244 19770 21303
rect 20108 21244 21598 21303
rect 22 21019 32 21172
rect 98 21019 108 21172
rect 214 21019 224 21172
rect 290 21019 300 21172
rect 406 21019 416 21172
rect 482 21019 492 21172
rect 598 21019 608 21172
rect 674 21019 684 21172
rect 790 21019 800 21172
rect 866 21019 876 21172
rect 982 21019 992 21172
rect 1058 21019 1068 21172
rect 1174 21019 1184 21172
rect 1250 21019 1260 21172
rect 1366 21019 1376 21172
rect 1442 21019 1452 21172
rect 1488 20959 1708 21206
rect 1850 21019 1860 21172
rect 1926 21019 1936 21172
rect 2042 21019 2052 21172
rect 2118 21019 2128 21172
rect 2234 21019 2244 21172
rect 2310 21019 2320 21172
rect 2426 21019 2436 21172
rect 2502 21019 2512 21172
rect 2618 21019 2628 21172
rect 2694 21019 2704 21172
rect 2810 21019 2820 21172
rect 2886 21019 2896 21172
rect 3002 21019 3012 21172
rect 3078 21019 3088 21172
rect 3194 21019 3204 21172
rect 3270 21019 3280 21172
rect 3316 20959 3536 21206
rect 3678 21019 3688 21172
rect 3754 21019 3764 21172
rect 3870 21019 3880 21172
rect 3946 21019 3956 21172
rect 4062 21019 4072 21172
rect 4138 21019 4148 21172
rect 4254 21019 4264 21172
rect 4330 21019 4340 21172
rect 4446 21019 4456 21172
rect 4522 21019 4532 21172
rect 4638 21019 4648 21172
rect 4714 21019 4724 21172
rect 4830 21019 4840 21172
rect 4906 21019 4916 21172
rect 5022 21019 5032 21172
rect 5098 21019 5108 21172
rect 5144 20959 5364 21206
rect 5506 21019 5516 21172
rect 5582 21019 5592 21172
rect 5698 21019 5708 21172
rect 5774 21019 5784 21172
rect 5890 21019 5900 21172
rect 5966 21019 5976 21172
rect 6082 21019 6092 21172
rect 6158 21019 6168 21172
rect 6274 21019 6284 21172
rect 6350 21019 6360 21172
rect 6466 21019 6476 21172
rect 6542 21019 6552 21172
rect 6658 21019 6668 21172
rect 6734 21019 6744 21172
rect 6850 21019 6860 21172
rect 6926 21019 6936 21172
rect 6972 20959 7192 21206
rect 7334 21019 7344 21172
rect 7410 21019 7420 21172
rect 7526 21019 7536 21172
rect 7602 21019 7612 21172
rect 7718 21019 7728 21172
rect 7794 21019 7804 21172
rect 7910 21019 7920 21172
rect 7986 21019 7996 21172
rect 8102 21019 8112 21172
rect 8178 21019 8188 21172
rect 8294 21019 8304 21172
rect 8370 21019 8380 21172
rect 8486 21019 8496 21172
rect 8562 21019 8572 21172
rect 8678 21019 8688 21172
rect 8754 21019 8764 21172
rect 8800 20959 9020 21206
rect 9162 21019 9172 21172
rect 9238 21019 9248 21172
rect 9354 21019 9364 21172
rect 9430 21019 9440 21172
rect 9546 21019 9556 21172
rect 9622 21019 9632 21172
rect 9738 21019 9748 21172
rect 9814 21019 9824 21172
rect 9930 21019 9940 21172
rect 10006 21019 10016 21172
rect 10122 21019 10132 21172
rect 10198 21019 10208 21172
rect 10314 21019 10324 21172
rect 10390 21019 10400 21172
rect 10506 21019 10516 21172
rect 10582 21019 10592 21172
rect 10628 20959 10848 21206
rect 10990 21019 11000 21172
rect 11066 21019 11076 21172
rect 11182 21019 11192 21172
rect 11258 21019 11268 21172
rect 11374 21019 11384 21172
rect 11450 21019 11460 21172
rect 11566 21019 11576 21172
rect 11642 21019 11652 21172
rect 11758 21019 11768 21172
rect 11834 21019 11844 21172
rect 11950 21019 11960 21172
rect 12026 21019 12036 21172
rect 12142 21019 12152 21172
rect 12218 21019 12228 21172
rect 12334 21019 12344 21172
rect 12410 21019 12420 21172
rect 12456 20959 12676 21206
rect 12818 21019 12828 21172
rect 12894 21019 12904 21172
rect 13010 21019 13020 21172
rect 13086 21019 13096 21172
rect 13202 21019 13212 21172
rect 13278 21019 13288 21172
rect 13394 21019 13404 21172
rect 13470 21019 13480 21172
rect 13586 21019 13596 21172
rect 13662 21019 13672 21172
rect 13778 21019 13788 21172
rect 13854 21019 13864 21172
rect 13970 21019 13980 21172
rect 14046 21019 14056 21172
rect 14162 21019 14172 21172
rect 14238 21019 14248 21172
rect 14284 20959 14504 21206
rect 14646 21019 14656 21172
rect 14722 21019 14732 21172
rect 14838 21019 14848 21172
rect 14914 21019 14924 21172
rect 15030 21019 15040 21172
rect 15106 21019 15116 21172
rect 15222 21019 15232 21172
rect 15298 21019 15308 21172
rect 15414 21019 15424 21172
rect 15490 21019 15500 21172
rect 15606 21019 15616 21172
rect 15682 21019 15692 21172
rect 15798 21019 15808 21172
rect 15874 21019 15884 21172
rect 15990 21019 16000 21172
rect 16066 21019 16076 21172
rect 16112 20959 16332 21206
rect 16474 21019 16484 21172
rect 16550 21019 16560 21172
rect 16666 21019 16676 21172
rect 16742 21019 16752 21172
rect 16858 21019 16868 21172
rect 16934 21019 16944 21172
rect 17050 21019 17060 21172
rect 17126 21019 17136 21172
rect 17242 21019 17252 21172
rect 17318 21019 17328 21172
rect 17434 21019 17444 21172
rect 17510 21019 17520 21172
rect 17626 21019 17636 21172
rect 17702 21019 17712 21172
rect 17818 21019 17828 21172
rect 17894 21019 17904 21172
rect 17940 20959 18160 21206
rect 18302 21019 18312 21172
rect 18378 21019 18388 21172
rect 18494 21019 18504 21172
rect 18570 21019 18580 21172
rect 18686 21019 18696 21172
rect 18762 21019 18772 21172
rect 18878 21019 18888 21172
rect 18954 21019 18964 21172
rect 19070 21019 19080 21172
rect 19146 21019 19156 21172
rect 19262 21019 19272 21172
rect 19338 21019 19348 21172
rect 19454 21019 19464 21172
rect 19530 21019 19540 21172
rect 19646 21019 19656 21172
rect 19722 21019 19732 21172
rect 19768 20959 19988 21206
rect 20130 21019 20140 21172
rect 20206 21019 20216 21172
rect 20322 21019 20332 21172
rect 20398 21019 20408 21172
rect 20514 21019 20524 21172
rect 20590 21019 20600 21172
rect 20706 21019 20716 21172
rect 20782 21019 20792 21172
rect 20898 21019 20908 21172
rect 20974 21019 20984 21172
rect 21090 21019 21100 21172
rect 21166 21019 21176 21172
rect 21282 21019 21292 21172
rect 21358 21019 21368 21172
rect 21474 21019 21484 21172
rect 21550 21019 21560 21172
rect 21596 20959 21816 21206
rect 118 20806 128 20959
rect 194 20806 204 20959
rect 310 20806 320 20959
rect 386 20806 396 20959
rect 502 20806 512 20959
rect 578 20806 588 20959
rect 694 20806 704 20959
rect 770 20806 780 20959
rect 886 20806 896 20959
rect 962 20806 972 20959
rect 1078 20806 1088 20959
rect 1154 20806 1164 20959
rect 1270 20806 1280 20959
rect 1346 20806 1356 20959
rect 1462 20806 1472 20959
rect 1528 20806 1708 20959
rect 1946 20806 1956 20959
rect 2022 20806 2032 20959
rect 2138 20806 2148 20959
rect 2214 20806 2224 20959
rect 2330 20806 2340 20959
rect 2406 20806 2416 20959
rect 2522 20806 2532 20959
rect 2598 20806 2608 20959
rect 2714 20806 2724 20959
rect 2790 20806 2800 20959
rect 2906 20806 2916 20959
rect 2982 20806 2992 20959
rect 3098 20806 3108 20959
rect 3174 20806 3184 20959
rect 3290 20806 3300 20959
rect 3356 20806 3536 20959
rect 3774 20806 3784 20959
rect 3850 20806 3860 20959
rect 3966 20806 3976 20959
rect 4042 20806 4052 20959
rect 4158 20806 4168 20959
rect 4234 20806 4244 20959
rect 4350 20806 4360 20959
rect 4426 20806 4436 20959
rect 4542 20806 4552 20959
rect 4618 20806 4628 20959
rect 4734 20806 4744 20959
rect 4810 20806 4820 20959
rect 4926 20806 4936 20959
rect 5002 20806 5012 20959
rect 5118 20806 5128 20959
rect 5184 20806 5364 20959
rect 5602 20806 5612 20959
rect 5678 20806 5688 20959
rect 5794 20806 5804 20959
rect 5870 20806 5880 20959
rect 5986 20806 5996 20959
rect 6062 20806 6072 20959
rect 6178 20806 6188 20959
rect 6254 20806 6264 20959
rect 6370 20806 6380 20959
rect 6446 20806 6456 20959
rect 6562 20806 6572 20959
rect 6638 20806 6648 20959
rect 6754 20806 6764 20959
rect 6830 20806 6840 20959
rect 6946 20806 6956 20959
rect 7012 20806 7192 20959
rect 7430 20806 7440 20959
rect 7506 20806 7516 20959
rect 7622 20806 7632 20959
rect 7698 20806 7708 20959
rect 7814 20806 7824 20959
rect 7890 20806 7900 20959
rect 8006 20806 8016 20959
rect 8082 20806 8092 20959
rect 8198 20806 8208 20959
rect 8274 20806 8284 20959
rect 8390 20806 8400 20959
rect 8466 20806 8476 20959
rect 8582 20806 8592 20959
rect 8658 20806 8668 20959
rect 8774 20806 8784 20959
rect 8840 20806 9020 20959
rect 9258 20806 9268 20959
rect 9334 20806 9344 20959
rect 9450 20806 9460 20959
rect 9526 20806 9536 20959
rect 9642 20806 9652 20959
rect 9718 20806 9728 20959
rect 9834 20806 9844 20959
rect 9910 20806 9920 20959
rect 10026 20806 10036 20959
rect 10102 20806 10112 20959
rect 10218 20806 10228 20959
rect 10294 20806 10304 20959
rect 10410 20806 10420 20959
rect 10486 20806 10496 20959
rect 10602 20806 10612 20959
rect 10668 20806 10848 20959
rect 11086 20806 11096 20959
rect 11162 20806 11172 20959
rect 11278 20806 11288 20959
rect 11354 20806 11364 20959
rect 11470 20806 11480 20959
rect 11546 20806 11556 20959
rect 11662 20806 11672 20959
rect 11738 20806 11748 20959
rect 11854 20806 11864 20959
rect 11930 20806 11940 20959
rect 12046 20806 12056 20959
rect 12122 20806 12132 20959
rect 12238 20806 12248 20959
rect 12314 20806 12324 20959
rect 12430 20806 12440 20959
rect 12496 20806 12676 20959
rect 12914 20806 12924 20959
rect 12990 20806 13000 20959
rect 13106 20806 13116 20959
rect 13182 20806 13192 20959
rect 13298 20806 13308 20959
rect 13374 20806 13384 20959
rect 13490 20806 13500 20959
rect 13566 20806 13576 20959
rect 13682 20806 13692 20959
rect 13758 20806 13768 20959
rect 13874 20806 13884 20959
rect 13950 20806 13960 20959
rect 14066 20806 14076 20959
rect 14142 20806 14152 20959
rect 14258 20806 14268 20959
rect 14324 20806 14504 20959
rect 14742 20806 14752 20959
rect 14818 20806 14828 20959
rect 14934 20806 14944 20959
rect 15010 20806 15020 20959
rect 15126 20806 15136 20959
rect 15202 20806 15212 20959
rect 15318 20806 15328 20959
rect 15394 20806 15404 20959
rect 15510 20806 15520 20959
rect 15586 20806 15596 20959
rect 15702 20806 15712 20959
rect 15778 20806 15788 20959
rect 15894 20806 15904 20959
rect 15970 20806 15980 20959
rect 16086 20806 16096 20959
rect 16152 20806 16332 20959
rect 16570 20806 16580 20959
rect 16646 20806 16656 20959
rect 16762 20806 16772 20959
rect 16838 20806 16848 20959
rect 16954 20806 16964 20959
rect 17030 20806 17040 20959
rect 17146 20806 17156 20959
rect 17222 20806 17232 20959
rect 17338 20806 17348 20959
rect 17414 20806 17424 20959
rect 17530 20806 17540 20959
rect 17606 20806 17616 20959
rect 17722 20806 17732 20959
rect 17798 20806 17808 20959
rect 17914 20806 17924 20959
rect 17980 20806 18160 20959
rect 18398 20806 18408 20959
rect 18474 20806 18484 20959
rect 18590 20806 18600 20959
rect 18666 20806 18676 20959
rect 18782 20806 18792 20959
rect 18858 20806 18868 20959
rect 18974 20806 18984 20959
rect 19050 20806 19060 20959
rect 19166 20806 19176 20959
rect 19242 20806 19252 20959
rect 19358 20806 19368 20959
rect 19434 20806 19444 20959
rect 19550 20806 19560 20959
rect 19626 20806 19636 20959
rect 19742 20806 19752 20959
rect 19808 20806 19988 20959
rect 20226 20806 20236 20959
rect 20302 20806 20312 20959
rect 20418 20806 20428 20959
rect 20494 20806 20504 20959
rect 20610 20806 20620 20959
rect 20686 20806 20696 20959
rect 20802 20806 20812 20959
rect 20878 20806 20888 20959
rect 20994 20806 21004 20959
rect 21070 20806 21080 20959
rect 21186 20806 21196 20959
rect 21262 20806 21272 20959
rect 21378 20806 21388 20959
rect 21454 20806 21464 20959
rect 21570 20806 21580 20959
rect 21636 20806 21816 20959
rect 0 20709 1490 20768
rect 1828 20709 3318 20768
rect 3656 20709 5146 20768
rect 5484 20709 6974 20768
rect 7312 20709 8802 20768
rect 9140 20709 10630 20768
rect 10968 20709 12458 20768
rect 12796 20709 14286 20768
rect 14624 20709 16114 20768
rect 16452 20709 17942 20768
rect 18280 20709 19770 20768
rect 20108 20709 21598 20768
rect 0 20530 1490 20589
rect 1828 20530 3318 20589
rect 3656 20530 5146 20589
rect 5484 20530 6974 20589
rect 7312 20530 8802 20589
rect 9140 20530 10630 20589
rect 10968 20530 12458 20589
rect 12796 20530 14286 20589
rect 14624 20530 16114 20589
rect 16452 20530 17942 20589
rect 18280 20530 19770 20589
rect 20108 20530 21598 20589
rect 22 20305 32 20458
rect 98 20305 108 20458
rect 214 20305 224 20458
rect 290 20305 300 20458
rect 406 20305 416 20458
rect 482 20305 492 20458
rect 598 20305 608 20458
rect 674 20305 684 20458
rect 790 20305 800 20458
rect 866 20305 876 20458
rect 982 20305 992 20458
rect 1058 20305 1068 20458
rect 1174 20305 1184 20458
rect 1250 20305 1260 20458
rect 1366 20305 1376 20458
rect 1442 20305 1452 20458
rect 1488 20245 1708 20492
rect 1850 20305 1860 20458
rect 1926 20305 1936 20458
rect 2042 20305 2052 20458
rect 2118 20305 2128 20458
rect 2234 20305 2244 20458
rect 2310 20305 2320 20458
rect 2426 20305 2436 20458
rect 2502 20305 2512 20458
rect 2618 20305 2628 20458
rect 2694 20305 2704 20458
rect 2810 20305 2820 20458
rect 2886 20305 2896 20458
rect 3002 20305 3012 20458
rect 3078 20305 3088 20458
rect 3194 20305 3204 20458
rect 3270 20305 3280 20458
rect 3316 20245 3536 20492
rect 3678 20305 3688 20458
rect 3754 20305 3764 20458
rect 3870 20305 3880 20458
rect 3946 20305 3956 20458
rect 4062 20305 4072 20458
rect 4138 20305 4148 20458
rect 4254 20305 4264 20458
rect 4330 20305 4340 20458
rect 4446 20305 4456 20458
rect 4522 20305 4532 20458
rect 4638 20305 4648 20458
rect 4714 20305 4724 20458
rect 4830 20305 4840 20458
rect 4906 20305 4916 20458
rect 5022 20305 5032 20458
rect 5098 20305 5108 20458
rect 5144 20245 5364 20492
rect 5506 20305 5516 20458
rect 5582 20305 5592 20458
rect 5698 20305 5708 20458
rect 5774 20305 5784 20458
rect 5890 20305 5900 20458
rect 5966 20305 5976 20458
rect 6082 20305 6092 20458
rect 6158 20305 6168 20458
rect 6274 20305 6284 20458
rect 6350 20305 6360 20458
rect 6466 20305 6476 20458
rect 6542 20305 6552 20458
rect 6658 20305 6668 20458
rect 6734 20305 6744 20458
rect 6850 20305 6860 20458
rect 6926 20305 6936 20458
rect 6972 20245 7192 20492
rect 7334 20305 7344 20458
rect 7410 20305 7420 20458
rect 7526 20305 7536 20458
rect 7602 20305 7612 20458
rect 7718 20305 7728 20458
rect 7794 20305 7804 20458
rect 7910 20305 7920 20458
rect 7986 20305 7996 20458
rect 8102 20305 8112 20458
rect 8178 20305 8188 20458
rect 8294 20305 8304 20458
rect 8370 20305 8380 20458
rect 8486 20305 8496 20458
rect 8562 20305 8572 20458
rect 8678 20305 8688 20458
rect 8754 20305 8764 20458
rect 8800 20245 9020 20492
rect 9162 20305 9172 20458
rect 9238 20305 9248 20458
rect 9354 20305 9364 20458
rect 9430 20305 9440 20458
rect 9546 20305 9556 20458
rect 9622 20305 9632 20458
rect 9738 20305 9748 20458
rect 9814 20305 9824 20458
rect 9930 20305 9940 20458
rect 10006 20305 10016 20458
rect 10122 20305 10132 20458
rect 10198 20305 10208 20458
rect 10314 20305 10324 20458
rect 10390 20305 10400 20458
rect 10506 20305 10516 20458
rect 10582 20305 10592 20458
rect 10628 20245 10848 20492
rect 10990 20305 11000 20458
rect 11066 20305 11076 20458
rect 11182 20305 11192 20458
rect 11258 20305 11268 20458
rect 11374 20305 11384 20458
rect 11450 20305 11460 20458
rect 11566 20305 11576 20458
rect 11642 20305 11652 20458
rect 11758 20305 11768 20458
rect 11834 20305 11844 20458
rect 11950 20305 11960 20458
rect 12026 20305 12036 20458
rect 12142 20305 12152 20458
rect 12218 20305 12228 20458
rect 12334 20305 12344 20458
rect 12410 20305 12420 20458
rect 12456 20245 12676 20492
rect 12818 20305 12828 20458
rect 12894 20305 12904 20458
rect 13010 20305 13020 20458
rect 13086 20305 13096 20458
rect 13202 20305 13212 20458
rect 13278 20305 13288 20458
rect 13394 20305 13404 20458
rect 13470 20305 13480 20458
rect 13586 20305 13596 20458
rect 13662 20305 13672 20458
rect 13778 20305 13788 20458
rect 13854 20305 13864 20458
rect 13970 20305 13980 20458
rect 14046 20305 14056 20458
rect 14162 20305 14172 20458
rect 14238 20305 14248 20458
rect 14284 20245 14504 20492
rect 14646 20305 14656 20458
rect 14722 20305 14732 20458
rect 14838 20305 14848 20458
rect 14914 20305 14924 20458
rect 15030 20305 15040 20458
rect 15106 20305 15116 20458
rect 15222 20305 15232 20458
rect 15298 20305 15308 20458
rect 15414 20305 15424 20458
rect 15490 20305 15500 20458
rect 15606 20305 15616 20458
rect 15682 20305 15692 20458
rect 15798 20305 15808 20458
rect 15874 20305 15884 20458
rect 15990 20305 16000 20458
rect 16066 20305 16076 20458
rect 16112 20245 16332 20492
rect 16474 20305 16484 20458
rect 16550 20305 16560 20458
rect 16666 20305 16676 20458
rect 16742 20305 16752 20458
rect 16858 20305 16868 20458
rect 16934 20305 16944 20458
rect 17050 20305 17060 20458
rect 17126 20305 17136 20458
rect 17242 20305 17252 20458
rect 17318 20305 17328 20458
rect 17434 20305 17444 20458
rect 17510 20305 17520 20458
rect 17626 20305 17636 20458
rect 17702 20305 17712 20458
rect 17818 20305 17828 20458
rect 17894 20305 17904 20458
rect 17940 20245 18160 20492
rect 18302 20305 18312 20458
rect 18378 20305 18388 20458
rect 18494 20305 18504 20458
rect 18570 20305 18580 20458
rect 18686 20305 18696 20458
rect 18762 20305 18772 20458
rect 18878 20305 18888 20458
rect 18954 20305 18964 20458
rect 19070 20305 19080 20458
rect 19146 20305 19156 20458
rect 19262 20305 19272 20458
rect 19338 20305 19348 20458
rect 19454 20305 19464 20458
rect 19530 20305 19540 20458
rect 19646 20305 19656 20458
rect 19722 20305 19732 20458
rect 19768 20245 19988 20492
rect 20130 20305 20140 20458
rect 20206 20305 20216 20458
rect 20322 20305 20332 20458
rect 20398 20305 20408 20458
rect 20514 20305 20524 20458
rect 20590 20305 20600 20458
rect 20706 20305 20716 20458
rect 20782 20305 20792 20458
rect 20898 20305 20908 20458
rect 20974 20305 20984 20458
rect 21090 20305 21100 20458
rect 21166 20305 21176 20458
rect 21282 20305 21292 20458
rect 21358 20305 21368 20458
rect 21474 20305 21484 20458
rect 21550 20305 21560 20458
rect 21596 20245 21816 20492
rect 118 20092 128 20245
rect 194 20092 204 20245
rect 310 20092 320 20245
rect 386 20092 396 20245
rect 502 20092 512 20245
rect 578 20092 588 20245
rect 694 20092 704 20245
rect 770 20092 780 20245
rect 886 20092 896 20245
rect 962 20092 972 20245
rect 1078 20092 1088 20245
rect 1154 20092 1164 20245
rect 1270 20092 1280 20245
rect 1346 20092 1356 20245
rect 1462 20092 1472 20245
rect 1528 20092 1708 20245
rect 1946 20092 1956 20245
rect 2022 20092 2032 20245
rect 2138 20092 2148 20245
rect 2214 20092 2224 20245
rect 2330 20092 2340 20245
rect 2406 20092 2416 20245
rect 2522 20092 2532 20245
rect 2598 20092 2608 20245
rect 2714 20092 2724 20245
rect 2790 20092 2800 20245
rect 2906 20092 2916 20245
rect 2982 20092 2992 20245
rect 3098 20092 3108 20245
rect 3174 20092 3184 20245
rect 3290 20092 3300 20245
rect 3356 20092 3536 20245
rect 3774 20092 3784 20245
rect 3850 20092 3860 20245
rect 3966 20092 3976 20245
rect 4042 20092 4052 20245
rect 4158 20092 4168 20245
rect 4234 20092 4244 20245
rect 4350 20092 4360 20245
rect 4426 20092 4436 20245
rect 4542 20092 4552 20245
rect 4618 20092 4628 20245
rect 4734 20092 4744 20245
rect 4810 20092 4820 20245
rect 4926 20092 4936 20245
rect 5002 20092 5012 20245
rect 5118 20092 5128 20245
rect 5184 20092 5364 20245
rect 5602 20092 5612 20245
rect 5678 20092 5688 20245
rect 5794 20092 5804 20245
rect 5870 20092 5880 20245
rect 5986 20092 5996 20245
rect 6062 20092 6072 20245
rect 6178 20092 6188 20245
rect 6254 20092 6264 20245
rect 6370 20092 6380 20245
rect 6446 20092 6456 20245
rect 6562 20092 6572 20245
rect 6638 20092 6648 20245
rect 6754 20092 6764 20245
rect 6830 20092 6840 20245
rect 6946 20092 6956 20245
rect 7012 20092 7192 20245
rect 7430 20092 7440 20245
rect 7506 20092 7516 20245
rect 7622 20092 7632 20245
rect 7698 20092 7708 20245
rect 7814 20092 7824 20245
rect 7890 20092 7900 20245
rect 8006 20092 8016 20245
rect 8082 20092 8092 20245
rect 8198 20092 8208 20245
rect 8274 20092 8284 20245
rect 8390 20092 8400 20245
rect 8466 20092 8476 20245
rect 8582 20092 8592 20245
rect 8658 20092 8668 20245
rect 8774 20092 8784 20245
rect 8840 20092 9020 20245
rect 9258 20092 9268 20245
rect 9334 20092 9344 20245
rect 9450 20092 9460 20245
rect 9526 20092 9536 20245
rect 9642 20092 9652 20245
rect 9718 20092 9728 20245
rect 9834 20092 9844 20245
rect 9910 20092 9920 20245
rect 10026 20092 10036 20245
rect 10102 20092 10112 20245
rect 10218 20092 10228 20245
rect 10294 20092 10304 20245
rect 10410 20092 10420 20245
rect 10486 20092 10496 20245
rect 10602 20092 10612 20245
rect 10668 20092 10848 20245
rect 11086 20092 11096 20245
rect 11162 20092 11172 20245
rect 11278 20092 11288 20245
rect 11354 20092 11364 20245
rect 11470 20092 11480 20245
rect 11546 20092 11556 20245
rect 11662 20092 11672 20245
rect 11738 20092 11748 20245
rect 11854 20092 11864 20245
rect 11930 20092 11940 20245
rect 12046 20092 12056 20245
rect 12122 20092 12132 20245
rect 12238 20092 12248 20245
rect 12314 20092 12324 20245
rect 12430 20092 12440 20245
rect 12496 20092 12676 20245
rect 12914 20092 12924 20245
rect 12990 20092 13000 20245
rect 13106 20092 13116 20245
rect 13182 20092 13192 20245
rect 13298 20092 13308 20245
rect 13374 20092 13384 20245
rect 13490 20092 13500 20245
rect 13566 20092 13576 20245
rect 13682 20092 13692 20245
rect 13758 20092 13768 20245
rect 13874 20092 13884 20245
rect 13950 20092 13960 20245
rect 14066 20092 14076 20245
rect 14142 20092 14152 20245
rect 14258 20092 14268 20245
rect 14324 20092 14504 20245
rect 14742 20092 14752 20245
rect 14818 20092 14828 20245
rect 14934 20092 14944 20245
rect 15010 20092 15020 20245
rect 15126 20092 15136 20245
rect 15202 20092 15212 20245
rect 15318 20092 15328 20245
rect 15394 20092 15404 20245
rect 15510 20092 15520 20245
rect 15586 20092 15596 20245
rect 15702 20092 15712 20245
rect 15778 20092 15788 20245
rect 15894 20092 15904 20245
rect 15970 20092 15980 20245
rect 16086 20092 16096 20245
rect 16152 20092 16332 20245
rect 16570 20092 16580 20245
rect 16646 20092 16656 20245
rect 16762 20092 16772 20245
rect 16838 20092 16848 20245
rect 16954 20092 16964 20245
rect 17030 20092 17040 20245
rect 17146 20092 17156 20245
rect 17222 20092 17232 20245
rect 17338 20092 17348 20245
rect 17414 20092 17424 20245
rect 17530 20092 17540 20245
rect 17606 20092 17616 20245
rect 17722 20092 17732 20245
rect 17798 20092 17808 20245
rect 17914 20092 17924 20245
rect 17980 20092 18160 20245
rect 18398 20092 18408 20245
rect 18474 20092 18484 20245
rect 18590 20092 18600 20245
rect 18666 20092 18676 20245
rect 18782 20092 18792 20245
rect 18858 20092 18868 20245
rect 18974 20092 18984 20245
rect 19050 20092 19060 20245
rect 19166 20092 19176 20245
rect 19242 20092 19252 20245
rect 19358 20092 19368 20245
rect 19434 20092 19444 20245
rect 19550 20092 19560 20245
rect 19626 20092 19636 20245
rect 19742 20092 19752 20245
rect 19808 20092 19988 20245
rect 20226 20092 20236 20245
rect 20302 20092 20312 20245
rect 20418 20092 20428 20245
rect 20494 20092 20504 20245
rect 20610 20092 20620 20245
rect 20686 20092 20696 20245
rect 20802 20092 20812 20245
rect 20878 20092 20888 20245
rect 20994 20092 21004 20245
rect 21070 20092 21080 20245
rect 21186 20092 21196 20245
rect 21262 20092 21272 20245
rect 21378 20092 21388 20245
rect 21454 20092 21464 20245
rect 21570 20092 21580 20245
rect 21636 20092 21816 20245
rect 0 19995 1490 20054
rect 1828 19995 3318 20054
rect 3656 19995 5146 20054
rect 5484 19995 6974 20054
rect 7312 19995 8802 20054
rect 9140 19995 10630 20054
rect 10968 19995 12458 20054
rect 12796 19995 14286 20054
rect 14624 19995 16114 20054
rect 16452 19995 17942 20054
rect 18280 19995 19770 20054
rect 20108 19995 21598 20054
rect 0 19816 1490 19875
rect 1828 19816 3318 19875
rect 3656 19816 5146 19875
rect 5484 19816 6974 19875
rect 7312 19816 8802 19875
rect 9140 19816 10630 19875
rect 10968 19816 12458 19875
rect 12796 19816 14286 19875
rect 14624 19816 16114 19875
rect 16452 19816 17942 19875
rect 18280 19816 19770 19875
rect 20108 19816 21598 19875
rect 22 19591 32 19744
rect 98 19591 108 19744
rect 214 19591 224 19744
rect 290 19591 300 19744
rect 406 19591 416 19744
rect 482 19591 492 19744
rect 598 19591 608 19744
rect 674 19591 684 19744
rect 790 19591 800 19744
rect 866 19591 876 19744
rect 982 19591 992 19744
rect 1058 19591 1068 19744
rect 1174 19591 1184 19744
rect 1250 19591 1260 19744
rect 1366 19591 1376 19744
rect 1442 19591 1452 19744
rect 1488 19531 1708 19778
rect 1850 19591 1860 19744
rect 1926 19591 1936 19744
rect 2042 19591 2052 19744
rect 2118 19591 2128 19744
rect 2234 19591 2244 19744
rect 2310 19591 2320 19744
rect 2426 19591 2436 19744
rect 2502 19591 2512 19744
rect 2618 19591 2628 19744
rect 2694 19591 2704 19744
rect 2810 19591 2820 19744
rect 2886 19591 2896 19744
rect 3002 19591 3012 19744
rect 3078 19591 3088 19744
rect 3194 19591 3204 19744
rect 3270 19591 3280 19744
rect 3316 19531 3536 19778
rect 3678 19591 3688 19744
rect 3754 19591 3764 19744
rect 3870 19591 3880 19744
rect 3946 19591 3956 19744
rect 4062 19591 4072 19744
rect 4138 19591 4148 19744
rect 4254 19591 4264 19744
rect 4330 19591 4340 19744
rect 4446 19591 4456 19744
rect 4522 19591 4532 19744
rect 4638 19591 4648 19744
rect 4714 19591 4724 19744
rect 4830 19591 4840 19744
rect 4906 19591 4916 19744
rect 5022 19591 5032 19744
rect 5098 19591 5108 19744
rect 5144 19531 5364 19778
rect 5506 19591 5516 19744
rect 5582 19591 5592 19744
rect 5698 19591 5708 19744
rect 5774 19591 5784 19744
rect 5890 19591 5900 19744
rect 5966 19591 5976 19744
rect 6082 19591 6092 19744
rect 6158 19591 6168 19744
rect 6274 19591 6284 19744
rect 6350 19591 6360 19744
rect 6466 19591 6476 19744
rect 6542 19591 6552 19744
rect 6658 19591 6668 19744
rect 6734 19591 6744 19744
rect 6850 19591 6860 19744
rect 6926 19591 6936 19744
rect 6972 19531 7192 19778
rect 7334 19591 7344 19744
rect 7410 19591 7420 19744
rect 7526 19591 7536 19744
rect 7602 19591 7612 19744
rect 7718 19591 7728 19744
rect 7794 19591 7804 19744
rect 7910 19591 7920 19744
rect 7986 19591 7996 19744
rect 8102 19591 8112 19744
rect 8178 19591 8188 19744
rect 8294 19591 8304 19744
rect 8370 19591 8380 19744
rect 8486 19591 8496 19744
rect 8562 19591 8572 19744
rect 8678 19591 8688 19744
rect 8754 19591 8764 19744
rect 8800 19531 9020 19778
rect 9162 19591 9172 19744
rect 9238 19591 9248 19744
rect 9354 19591 9364 19744
rect 9430 19591 9440 19744
rect 9546 19591 9556 19744
rect 9622 19591 9632 19744
rect 9738 19591 9748 19744
rect 9814 19591 9824 19744
rect 9930 19591 9940 19744
rect 10006 19591 10016 19744
rect 10122 19591 10132 19744
rect 10198 19591 10208 19744
rect 10314 19591 10324 19744
rect 10390 19591 10400 19744
rect 10506 19591 10516 19744
rect 10582 19591 10592 19744
rect 10628 19531 10848 19778
rect 10990 19591 11000 19744
rect 11066 19591 11076 19744
rect 11182 19591 11192 19744
rect 11258 19591 11268 19744
rect 11374 19591 11384 19744
rect 11450 19591 11460 19744
rect 11566 19591 11576 19744
rect 11642 19591 11652 19744
rect 11758 19591 11768 19744
rect 11834 19591 11844 19744
rect 11950 19591 11960 19744
rect 12026 19591 12036 19744
rect 12142 19591 12152 19744
rect 12218 19591 12228 19744
rect 12334 19591 12344 19744
rect 12410 19591 12420 19744
rect 12456 19531 12676 19778
rect 12818 19591 12828 19744
rect 12894 19591 12904 19744
rect 13010 19591 13020 19744
rect 13086 19591 13096 19744
rect 13202 19591 13212 19744
rect 13278 19591 13288 19744
rect 13394 19591 13404 19744
rect 13470 19591 13480 19744
rect 13586 19591 13596 19744
rect 13662 19591 13672 19744
rect 13778 19591 13788 19744
rect 13854 19591 13864 19744
rect 13970 19591 13980 19744
rect 14046 19591 14056 19744
rect 14162 19591 14172 19744
rect 14238 19591 14248 19744
rect 14284 19531 14504 19778
rect 14646 19591 14656 19744
rect 14722 19591 14732 19744
rect 14838 19591 14848 19744
rect 14914 19591 14924 19744
rect 15030 19591 15040 19744
rect 15106 19591 15116 19744
rect 15222 19591 15232 19744
rect 15298 19591 15308 19744
rect 15414 19591 15424 19744
rect 15490 19591 15500 19744
rect 15606 19591 15616 19744
rect 15682 19591 15692 19744
rect 15798 19591 15808 19744
rect 15874 19591 15884 19744
rect 15990 19591 16000 19744
rect 16066 19591 16076 19744
rect 16112 19531 16332 19778
rect 16474 19591 16484 19744
rect 16550 19591 16560 19744
rect 16666 19591 16676 19744
rect 16742 19591 16752 19744
rect 16858 19591 16868 19744
rect 16934 19591 16944 19744
rect 17050 19591 17060 19744
rect 17126 19591 17136 19744
rect 17242 19591 17252 19744
rect 17318 19591 17328 19744
rect 17434 19591 17444 19744
rect 17510 19591 17520 19744
rect 17626 19591 17636 19744
rect 17702 19591 17712 19744
rect 17818 19591 17828 19744
rect 17894 19591 17904 19744
rect 17940 19531 18160 19778
rect 18302 19591 18312 19744
rect 18378 19591 18388 19744
rect 18494 19591 18504 19744
rect 18570 19591 18580 19744
rect 18686 19591 18696 19744
rect 18762 19591 18772 19744
rect 18878 19591 18888 19744
rect 18954 19591 18964 19744
rect 19070 19591 19080 19744
rect 19146 19591 19156 19744
rect 19262 19591 19272 19744
rect 19338 19591 19348 19744
rect 19454 19591 19464 19744
rect 19530 19591 19540 19744
rect 19646 19591 19656 19744
rect 19722 19591 19732 19744
rect 19768 19531 19988 19778
rect 20130 19591 20140 19744
rect 20206 19591 20216 19744
rect 20322 19591 20332 19744
rect 20398 19591 20408 19744
rect 20514 19591 20524 19744
rect 20590 19591 20600 19744
rect 20706 19591 20716 19744
rect 20782 19591 20792 19744
rect 20898 19591 20908 19744
rect 20974 19591 20984 19744
rect 21090 19591 21100 19744
rect 21166 19591 21176 19744
rect 21282 19591 21292 19744
rect 21358 19591 21368 19744
rect 21474 19591 21484 19744
rect 21550 19591 21560 19744
rect 21596 19531 21816 19778
rect 118 19378 128 19531
rect 194 19378 204 19531
rect 310 19378 320 19531
rect 386 19378 396 19531
rect 502 19378 512 19531
rect 578 19378 588 19531
rect 694 19378 704 19531
rect 770 19378 780 19531
rect 886 19378 896 19531
rect 962 19378 972 19531
rect 1078 19378 1088 19531
rect 1154 19378 1164 19531
rect 1270 19378 1280 19531
rect 1346 19378 1356 19531
rect 1462 19378 1472 19531
rect 1528 19378 1708 19531
rect 1946 19378 1956 19531
rect 2022 19378 2032 19531
rect 2138 19378 2148 19531
rect 2214 19378 2224 19531
rect 2330 19378 2340 19531
rect 2406 19378 2416 19531
rect 2522 19378 2532 19531
rect 2598 19378 2608 19531
rect 2714 19378 2724 19531
rect 2790 19378 2800 19531
rect 2906 19378 2916 19531
rect 2982 19378 2992 19531
rect 3098 19378 3108 19531
rect 3174 19378 3184 19531
rect 3290 19378 3300 19531
rect 3356 19378 3536 19531
rect 3774 19378 3784 19531
rect 3850 19378 3860 19531
rect 3966 19378 3976 19531
rect 4042 19378 4052 19531
rect 4158 19378 4168 19531
rect 4234 19378 4244 19531
rect 4350 19378 4360 19531
rect 4426 19378 4436 19531
rect 4542 19378 4552 19531
rect 4618 19378 4628 19531
rect 4734 19378 4744 19531
rect 4810 19378 4820 19531
rect 4926 19378 4936 19531
rect 5002 19378 5012 19531
rect 5118 19378 5128 19531
rect 5184 19378 5364 19531
rect 5602 19378 5612 19531
rect 5678 19378 5688 19531
rect 5794 19378 5804 19531
rect 5870 19378 5880 19531
rect 5986 19378 5996 19531
rect 6062 19378 6072 19531
rect 6178 19378 6188 19531
rect 6254 19378 6264 19531
rect 6370 19378 6380 19531
rect 6446 19378 6456 19531
rect 6562 19378 6572 19531
rect 6638 19378 6648 19531
rect 6754 19378 6764 19531
rect 6830 19378 6840 19531
rect 6946 19378 6956 19531
rect 7012 19378 7192 19531
rect 7430 19378 7440 19531
rect 7506 19378 7516 19531
rect 7622 19378 7632 19531
rect 7698 19378 7708 19531
rect 7814 19378 7824 19531
rect 7890 19378 7900 19531
rect 8006 19378 8016 19531
rect 8082 19378 8092 19531
rect 8198 19378 8208 19531
rect 8274 19378 8284 19531
rect 8390 19378 8400 19531
rect 8466 19378 8476 19531
rect 8582 19378 8592 19531
rect 8658 19378 8668 19531
rect 8774 19378 8784 19531
rect 8840 19378 9020 19531
rect 9258 19378 9268 19531
rect 9334 19378 9344 19531
rect 9450 19378 9460 19531
rect 9526 19378 9536 19531
rect 9642 19378 9652 19531
rect 9718 19378 9728 19531
rect 9834 19378 9844 19531
rect 9910 19378 9920 19531
rect 10026 19378 10036 19531
rect 10102 19378 10112 19531
rect 10218 19378 10228 19531
rect 10294 19378 10304 19531
rect 10410 19378 10420 19531
rect 10486 19378 10496 19531
rect 10602 19378 10612 19531
rect 10668 19378 10848 19531
rect 11086 19378 11096 19531
rect 11162 19378 11172 19531
rect 11278 19378 11288 19531
rect 11354 19378 11364 19531
rect 11470 19378 11480 19531
rect 11546 19378 11556 19531
rect 11662 19378 11672 19531
rect 11738 19378 11748 19531
rect 11854 19378 11864 19531
rect 11930 19378 11940 19531
rect 12046 19378 12056 19531
rect 12122 19378 12132 19531
rect 12238 19378 12248 19531
rect 12314 19378 12324 19531
rect 12430 19378 12440 19531
rect 12496 19378 12676 19531
rect 12914 19378 12924 19531
rect 12990 19378 13000 19531
rect 13106 19378 13116 19531
rect 13182 19378 13192 19531
rect 13298 19378 13308 19531
rect 13374 19378 13384 19531
rect 13490 19378 13500 19531
rect 13566 19378 13576 19531
rect 13682 19378 13692 19531
rect 13758 19378 13768 19531
rect 13874 19378 13884 19531
rect 13950 19378 13960 19531
rect 14066 19378 14076 19531
rect 14142 19378 14152 19531
rect 14258 19378 14268 19531
rect 14324 19378 14504 19531
rect 14742 19378 14752 19531
rect 14818 19378 14828 19531
rect 14934 19378 14944 19531
rect 15010 19378 15020 19531
rect 15126 19378 15136 19531
rect 15202 19378 15212 19531
rect 15318 19378 15328 19531
rect 15394 19378 15404 19531
rect 15510 19378 15520 19531
rect 15586 19378 15596 19531
rect 15702 19378 15712 19531
rect 15778 19378 15788 19531
rect 15894 19378 15904 19531
rect 15970 19378 15980 19531
rect 16086 19378 16096 19531
rect 16152 19378 16332 19531
rect 16570 19378 16580 19531
rect 16646 19378 16656 19531
rect 16762 19378 16772 19531
rect 16838 19378 16848 19531
rect 16954 19378 16964 19531
rect 17030 19378 17040 19531
rect 17146 19378 17156 19531
rect 17222 19378 17232 19531
rect 17338 19378 17348 19531
rect 17414 19378 17424 19531
rect 17530 19378 17540 19531
rect 17606 19378 17616 19531
rect 17722 19378 17732 19531
rect 17798 19378 17808 19531
rect 17914 19378 17924 19531
rect 17980 19378 18160 19531
rect 18398 19378 18408 19531
rect 18474 19378 18484 19531
rect 18590 19378 18600 19531
rect 18666 19378 18676 19531
rect 18782 19378 18792 19531
rect 18858 19378 18868 19531
rect 18974 19378 18984 19531
rect 19050 19378 19060 19531
rect 19166 19378 19176 19531
rect 19242 19378 19252 19531
rect 19358 19378 19368 19531
rect 19434 19378 19444 19531
rect 19550 19378 19560 19531
rect 19626 19378 19636 19531
rect 19742 19378 19752 19531
rect 19808 19378 19988 19531
rect 20226 19378 20236 19531
rect 20302 19378 20312 19531
rect 20418 19378 20428 19531
rect 20494 19378 20504 19531
rect 20610 19378 20620 19531
rect 20686 19378 20696 19531
rect 20802 19378 20812 19531
rect 20878 19378 20888 19531
rect 20994 19378 21004 19531
rect 21070 19378 21080 19531
rect 21186 19378 21196 19531
rect 21262 19378 21272 19531
rect 21378 19378 21388 19531
rect 21454 19378 21464 19531
rect 21570 19378 21580 19531
rect 21636 19378 21816 19531
rect 0 19281 1490 19340
rect 1828 19281 3318 19340
rect 3656 19281 5146 19340
rect 5484 19281 6974 19340
rect 7312 19281 8802 19340
rect 9140 19281 10630 19340
rect 10968 19281 12458 19340
rect 12796 19281 14286 19340
rect 14624 19281 16114 19340
rect 16452 19281 17942 19340
rect 18280 19281 19770 19340
rect 20108 19281 21598 19340
rect 0 19102 1490 19161
rect 1828 19102 3318 19161
rect 3656 19102 5146 19161
rect 5484 19102 6974 19161
rect 7312 19102 8802 19161
rect 9140 19102 10630 19161
rect 10968 19102 12458 19161
rect 12796 19102 14286 19161
rect 14624 19102 16114 19161
rect 16452 19102 17942 19161
rect 18280 19102 19770 19161
rect 20108 19102 21598 19161
rect 22 18877 32 19030
rect 98 18877 108 19030
rect 214 18877 224 19030
rect 290 18877 300 19030
rect 406 18877 416 19030
rect 482 18877 492 19030
rect 598 18877 608 19030
rect 674 18877 684 19030
rect 790 18877 800 19030
rect 866 18877 876 19030
rect 982 18877 992 19030
rect 1058 18877 1068 19030
rect 1174 18877 1184 19030
rect 1250 18877 1260 19030
rect 1366 18877 1376 19030
rect 1442 18877 1452 19030
rect 1488 18817 1708 19064
rect 1850 18877 1860 19030
rect 1926 18877 1936 19030
rect 2042 18877 2052 19030
rect 2118 18877 2128 19030
rect 2234 18877 2244 19030
rect 2310 18877 2320 19030
rect 2426 18877 2436 19030
rect 2502 18877 2512 19030
rect 2618 18877 2628 19030
rect 2694 18877 2704 19030
rect 2810 18877 2820 19030
rect 2886 18877 2896 19030
rect 3002 18877 3012 19030
rect 3078 18877 3088 19030
rect 3194 18877 3204 19030
rect 3270 18877 3280 19030
rect 3316 18817 3536 19064
rect 3678 18877 3688 19030
rect 3754 18877 3764 19030
rect 3870 18877 3880 19030
rect 3946 18877 3956 19030
rect 4062 18877 4072 19030
rect 4138 18877 4148 19030
rect 4254 18877 4264 19030
rect 4330 18877 4340 19030
rect 4446 18877 4456 19030
rect 4522 18877 4532 19030
rect 4638 18877 4648 19030
rect 4714 18877 4724 19030
rect 4830 18877 4840 19030
rect 4906 18877 4916 19030
rect 5022 18877 5032 19030
rect 5098 18877 5108 19030
rect 5144 18817 5364 19064
rect 5506 18877 5516 19030
rect 5582 18877 5592 19030
rect 5698 18877 5708 19030
rect 5774 18877 5784 19030
rect 5890 18877 5900 19030
rect 5966 18877 5976 19030
rect 6082 18877 6092 19030
rect 6158 18877 6168 19030
rect 6274 18877 6284 19030
rect 6350 18877 6360 19030
rect 6466 18877 6476 19030
rect 6542 18877 6552 19030
rect 6658 18877 6668 19030
rect 6734 18877 6744 19030
rect 6850 18877 6860 19030
rect 6926 18877 6936 19030
rect 6972 18817 7192 19064
rect 7334 18877 7344 19030
rect 7410 18877 7420 19030
rect 7526 18877 7536 19030
rect 7602 18877 7612 19030
rect 7718 18877 7728 19030
rect 7794 18877 7804 19030
rect 7910 18877 7920 19030
rect 7986 18877 7996 19030
rect 8102 18877 8112 19030
rect 8178 18877 8188 19030
rect 8294 18877 8304 19030
rect 8370 18877 8380 19030
rect 8486 18877 8496 19030
rect 8562 18877 8572 19030
rect 8678 18877 8688 19030
rect 8754 18877 8764 19030
rect 8800 18817 9020 19064
rect 9162 18877 9172 19030
rect 9238 18877 9248 19030
rect 9354 18877 9364 19030
rect 9430 18877 9440 19030
rect 9546 18877 9556 19030
rect 9622 18877 9632 19030
rect 9738 18877 9748 19030
rect 9814 18877 9824 19030
rect 9930 18877 9940 19030
rect 10006 18877 10016 19030
rect 10122 18877 10132 19030
rect 10198 18877 10208 19030
rect 10314 18877 10324 19030
rect 10390 18877 10400 19030
rect 10506 18877 10516 19030
rect 10582 18877 10592 19030
rect 10628 18817 10848 19064
rect 10990 18877 11000 19030
rect 11066 18877 11076 19030
rect 11182 18877 11192 19030
rect 11258 18877 11268 19030
rect 11374 18877 11384 19030
rect 11450 18877 11460 19030
rect 11566 18877 11576 19030
rect 11642 18877 11652 19030
rect 11758 18877 11768 19030
rect 11834 18877 11844 19030
rect 11950 18877 11960 19030
rect 12026 18877 12036 19030
rect 12142 18877 12152 19030
rect 12218 18877 12228 19030
rect 12334 18877 12344 19030
rect 12410 18877 12420 19030
rect 12456 18817 12676 19064
rect 12818 18877 12828 19030
rect 12894 18877 12904 19030
rect 13010 18877 13020 19030
rect 13086 18877 13096 19030
rect 13202 18877 13212 19030
rect 13278 18877 13288 19030
rect 13394 18877 13404 19030
rect 13470 18877 13480 19030
rect 13586 18877 13596 19030
rect 13662 18877 13672 19030
rect 13778 18877 13788 19030
rect 13854 18877 13864 19030
rect 13970 18877 13980 19030
rect 14046 18877 14056 19030
rect 14162 18877 14172 19030
rect 14238 18877 14248 19030
rect 14284 18817 14504 19064
rect 14646 18877 14656 19030
rect 14722 18877 14732 19030
rect 14838 18877 14848 19030
rect 14914 18877 14924 19030
rect 15030 18877 15040 19030
rect 15106 18877 15116 19030
rect 15222 18877 15232 19030
rect 15298 18877 15308 19030
rect 15414 18877 15424 19030
rect 15490 18877 15500 19030
rect 15606 18877 15616 19030
rect 15682 18877 15692 19030
rect 15798 18877 15808 19030
rect 15874 18877 15884 19030
rect 15990 18877 16000 19030
rect 16066 18877 16076 19030
rect 16112 18817 16332 19064
rect 16474 18877 16484 19030
rect 16550 18877 16560 19030
rect 16666 18877 16676 19030
rect 16742 18877 16752 19030
rect 16858 18877 16868 19030
rect 16934 18877 16944 19030
rect 17050 18877 17060 19030
rect 17126 18877 17136 19030
rect 17242 18877 17252 19030
rect 17318 18877 17328 19030
rect 17434 18877 17444 19030
rect 17510 18877 17520 19030
rect 17626 18877 17636 19030
rect 17702 18877 17712 19030
rect 17818 18877 17828 19030
rect 17894 18877 17904 19030
rect 17940 18817 18160 19064
rect 18302 18877 18312 19030
rect 18378 18877 18388 19030
rect 18494 18877 18504 19030
rect 18570 18877 18580 19030
rect 18686 18877 18696 19030
rect 18762 18877 18772 19030
rect 18878 18877 18888 19030
rect 18954 18877 18964 19030
rect 19070 18877 19080 19030
rect 19146 18877 19156 19030
rect 19262 18877 19272 19030
rect 19338 18877 19348 19030
rect 19454 18877 19464 19030
rect 19530 18877 19540 19030
rect 19646 18877 19656 19030
rect 19722 18877 19732 19030
rect 19768 18817 19988 19064
rect 20130 18877 20140 19030
rect 20206 18877 20216 19030
rect 20322 18877 20332 19030
rect 20398 18877 20408 19030
rect 20514 18877 20524 19030
rect 20590 18877 20600 19030
rect 20706 18877 20716 19030
rect 20782 18877 20792 19030
rect 20898 18877 20908 19030
rect 20974 18877 20984 19030
rect 21090 18877 21100 19030
rect 21166 18877 21176 19030
rect 21282 18877 21292 19030
rect 21358 18877 21368 19030
rect 21474 18877 21484 19030
rect 21550 18877 21560 19030
rect 21596 18817 21816 19064
rect 118 18664 128 18817
rect 194 18664 204 18817
rect 310 18664 320 18817
rect 386 18664 396 18817
rect 502 18664 512 18817
rect 578 18664 588 18817
rect 694 18664 704 18817
rect 770 18664 780 18817
rect 886 18664 896 18817
rect 962 18664 972 18817
rect 1078 18664 1088 18817
rect 1154 18664 1164 18817
rect 1270 18664 1280 18817
rect 1346 18664 1356 18817
rect 1462 18664 1472 18817
rect 1528 18664 1708 18817
rect 1946 18664 1956 18817
rect 2022 18664 2032 18817
rect 2138 18664 2148 18817
rect 2214 18664 2224 18817
rect 2330 18664 2340 18817
rect 2406 18664 2416 18817
rect 2522 18664 2532 18817
rect 2598 18664 2608 18817
rect 2714 18664 2724 18817
rect 2790 18664 2800 18817
rect 2906 18664 2916 18817
rect 2982 18664 2992 18817
rect 3098 18664 3108 18817
rect 3174 18664 3184 18817
rect 3290 18664 3300 18817
rect 3356 18664 3536 18817
rect 3774 18664 3784 18817
rect 3850 18664 3860 18817
rect 3966 18664 3976 18817
rect 4042 18664 4052 18817
rect 4158 18664 4168 18817
rect 4234 18664 4244 18817
rect 4350 18664 4360 18817
rect 4426 18664 4436 18817
rect 4542 18664 4552 18817
rect 4618 18664 4628 18817
rect 4734 18664 4744 18817
rect 4810 18664 4820 18817
rect 4926 18664 4936 18817
rect 5002 18664 5012 18817
rect 5118 18664 5128 18817
rect 5184 18664 5364 18817
rect 5602 18664 5612 18817
rect 5678 18664 5688 18817
rect 5794 18664 5804 18817
rect 5870 18664 5880 18817
rect 5986 18664 5996 18817
rect 6062 18664 6072 18817
rect 6178 18664 6188 18817
rect 6254 18664 6264 18817
rect 6370 18664 6380 18817
rect 6446 18664 6456 18817
rect 6562 18664 6572 18817
rect 6638 18664 6648 18817
rect 6754 18664 6764 18817
rect 6830 18664 6840 18817
rect 6946 18664 6956 18817
rect 7012 18664 7192 18817
rect 7430 18664 7440 18817
rect 7506 18664 7516 18817
rect 7622 18664 7632 18817
rect 7698 18664 7708 18817
rect 7814 18664 7824 18817
rect 7890 18664 7900 18817
rect 8006 18664 8016 18817
rect 8082 18664 8092 18817
rect 8198 18664 8208 18817
rect 8274 18664 8284 18817
rect 8390 18664 8400 18817
rect 8466 18664 8476 18817
rect 8582 18664 8592 18817
rect 8658 18664 8668 18817
rect 8774 18664 8784 18817
rect 8840 18664 9020 18817
rect 9258 18664 9268 18817
rect 9334 18664 9344 18817
rect 9450 18664 9460 18817
rect 9526 18664 9536 18817
rect 9642 18664 9652 18817
rect 9718 18664 9728 18817
rect 9834 18664 9844 18817
rect 9910 18664 9920 18817
rect 10026 18664 10036 18817
rect 10102 18664 10112 18817
rect 10218 18664 10228 18817
rect 10294 18664 10304 18817
rect 10410 18664 10420 18817
rect 10486 18664 10496 18817
rect 10602 18664 10612 18817
rect 10668 18664 10848 18817
rect 11086 18664 11096 18817
rect 11162 18664 11172 18817
rect 11278 18664 11288 18817
rect 11354 18664 11364 18817
rect 11470 18664 11480 18817
rect 11546 18664 11556 18817
rect 11662 18664 11672 18817
rect 11738 18664 11748 18817
rect 11854 18664 11864 18817
rect 11930 18664 11940 18817
rect 12046 18664 12056 18817
rect 12122 18664 12132 18817
rect 12238 18664 12248 18817
rect 12314 18664 12324 18817
rect 12430 18664 12440 18817
rect 12496 18664 12676 18817
rect 12914 18664 12924 18817
rect 12990 18664 13000 18817
rect 13106 18664 13116 18817
rect 13182 18664 13192 18817
rect 13298 18664 13308 18817
rect 13374 18664 13384 18817
rect 13490 18664 13500 18817
rect 13566 18664 13576 18817
rect 13682 18664 13692 18817
rect 13758 18664 13768 18817
rect 13874 18664 13884 18817
rect 13950 18664 13960 18817
rect 14066 18664 14076 18817
rect 14142 18664 14152 18817
rect 14258 18664 14268 18817
rect 14324 18664 14504 18817
rect 14742 18664 14752 18817
rect 14818 18664 14828 18817
rect 14934 18664 14944 18817
rect 15010 18664 15020 18817
rect 15126 18664 15136 18817
rect 15202 18664 15212 18817
rect 15318 18664 15328 18817
rect 15394 18664 15404 18817
rect 15510 18664 15520 18817
rect 15586 18664 15596 18817
rect 15702 18664 15712 18817
rect 15778 18664 15788 18817
rect 15894 18664 15904 18817
rect 15970 18664 15980 18817
rect 16086 18664 16096 18817
rect 16152 18664 16332 18817
rect 16570 18664 16580 18817
rect 16646 18664 16656 18817
rect 16762 18664 16772 18817
rect 16838 18664 16848 18817
rect 16954 18664 16964 18817
rect 17030 18664 17040 18817
rect 17146 18664 17156 18817
rect 17222 18664 17232 18817
rect 17338 18664 17348 18817
rect 17414 18664 17424 18817
rect 17530 18664 17540 18817
rect 17606 18664 17616 18817
rect 17722 18664 17732 18817
rect 17798 18664 17808 18817
rect 17914 18664 17924 18817
rect 17980 18664 18160 18817
rect 18398 18664 18408 18817
rect 18474 18664 18484 18817
rect 18590 18664 18600 18817
rect 18666 18664 18676 18817
rect 18782 18664 18792 18817
rect 18858 18664 18868 18817
rect 18974 18664 18984 18817
rect 19050 18664 19060 18817
rect 19166 18664 19176 18817
rect 19242 18664 19252 18817
rect 19358 18664 19368 18817
rect 19434 18664 19444 18817
rect 19550 18664 19560 18817
rect 19626 18664 19636 18817
rect 19742 18664 19752 18817
rect 19808 18664 19988 18817
rect 20226 18664 20236 18817
rect 20302 18664 20312 18817
rect 20418 18664 20428 18817
rect 20494 18664 20504 18817
rect 20610 18664 20620 18817
rect 20686 18664 20696 18817
rect 20802 18664 20812 18817
rect 20878 18664 20888 18817
rect 20994 18664 21004 18817
rect 21070 18664 21080 18817
rect 21186 18664 21196 18817
rect 21262 18664 21272 18817
rect 21378 18664 21388 18817
rect 21454 18664 21464 18817
rect 21570 18664 21580 18817
rect 21636 18664 21816 18817
rect 0 18567 1490 18626
rect 1828 18567 3318 18626
rect 3656 18567 5146 18626
rect 5484 18567 6974 18626
rect 7312 18567 8802 18626
rect 9140 18567 10630 18626
rect 10968 18567 12458 18626
rect 12796 18567 14286 18626
rect 14624 18567 16114 18626
rect 16452 18567 17942 18626
rect 18280 18567 19770 18626
rect 20108 18567 21598 18626
rect 0 18388 1490 18447
rect 1828 18388 3318 18447
rect 3656 18388 5146 18447
rect 5484 18388 6974 18447
rect 7312 18388 8802 18447
rect 9140 18388 10630 18447
rect 10968 18388 12458 18447
rect 12796 18388 14286 18447
rect 14624 18388 16114 18447
rect 16452 18388 17942 18447
rect 18280 18388 19770 18447
rect 20108 18388 21598 18447
rect 22 18163 32 18316
rect 98 18163 108 18316
rect 214 18163 224 18316
rect 290 18163 300 18316
rect 406 18163 416 18316
rect 482 18163 492 18316
rect 598 18163 608 18316
rect 674 18163 684 18316
rect 790 18163 800 18316
rect 866 18163 876 18316
rect 982 18163 992 18316
rect 1058 18163 1068 18316
rect 1174 18163 1184 18316
rect 1250 18163 1260 18316
rect 1366 18163 1376 18316
rect 1442 18163 1452 18316
rect 1488 18103 1708 18350
rect 1850 18163 1860 18316
rect 1926 18163 1936 18316
rect 2042 18163 2052 18316
rect 2118 18163 2128 18316
rect 2234 18163 2244 18316
rect 2310 18163 2320 18316
rect 2426 18163 2436 18316
rect 2502 18163 2512 18316
rect 2618 18163 2628 18316
rect 2694 18163 2704 18316
rect 2810 18163 2820 18316
rect 2886 18163 2896 18316
rect 3002 18163 3012 18316
rect 3078 18163 3088 18316
rect 3194 18163 3204 18316
rect 3270 18163 3280 18316
rect 3316 18103 3536 18350
rect 3678 18163 3688 18316
rect 3754 18163 3764 18316
rect 3870 18163 3880 18316
rect 3946 18163 3956 18316
rect 4062 18163 4072 18316
rect 4138 18163 4148 18316
rect 4254 18163 4264 18316
rect 4330 18163 4340 18316
rect 4446 18163 4456 18316
rect 4522 18163 4532 18316
rect 4638 18163 4648 18316
rect 4714 18163 4724 18316
rect 4830 18163 4840 18316
rect 4906 18163 4916 18316
rect 5022 18163 5032 18316
rect 5098 18163 5108 18316
rect 5144 18103 5364 18350
rect 5506 18163 5516 18316
rect 5582 18163 5592 18316
rect 5698 18163 5708 18316
rect 5774 18163 5784 18316
rect 5890 18163 5900 18316
rect 5966 18163 5976 18316
rect 6082 18163 6092 18316
rect 6158 18163 6168 18316
rect 6274 18163 6284 18316
rect 6350 18163 6360 18316
rect 6466 18163 6476 18316
rect 6542 18163 6552 18316
rect 6658 18163 6668 18316
rect 6734 18163 6744 18316
rect 6850 18163 6860 18316
rect 6926 18163 6936 18316
rect 6972 18103 7192 18350
rect 7334 18163 7344 18316
rect 7410 18163 7420 18316
rect 7526 18163 7536 18316
rect 7602 18163 7612 18316
rect 7718 18163 7728 18316
rect 7794 18163 7804 18316
rect 7910 18163 7920 18316
rect 7986 18163 7996 18316
rect 8102 18163 8112 18316
rect 8178 18163 8188 18316
rect 8294 18163 8304 18316
rect 8370 18163 8380 18316
rect 8486 18163 8496 18316
rect 8562 18163 8572 18316
rect 8678 18163 8688 18316
rect 8754 18163 8764 18316
rect 8800 18103 9020 18350
rect 9162 18163 9172 18316
rect 9238 18163 9248 18316
rect 9354 18163 9364 18316
rect 9430 18163 9440 18316
rect 9546 18163 9556 18316
rect 9622 18163 9632 18316
rect 9738 18163 9748 18316
rect 9814 18163 9824 18316
rect 9930 18163 9940 18316
rect 10006 18163 10016 18316
rect 10122 18163 10132 18316
rect 10198 18163 10208 18316
rect 10314 18163 10324 18316
rect 10390 18163 10400 18316
rect 10506 18163 10516 18316
rect 10582 18163 10592 18316
rect 10628 18103 10848 18350
rect 10990 18163 11000 18316
rect 11066 18163 11076 18316
rect 11182 18163 11192 18316
rect 11258 18163 11268 18316
rect 11374 18163 11384 18316
rect 11450 18163 11460 18316
rect 11566 18163 11576 18316
rect 11642 18163 11652 18316
rect 11758 18163 11768 18316
rect 11834 18163 11844 18316
rect 11950 18163 11960 18316
rect 12026 18163 12036 18316
rect 12142 18163 12152 18316
rect 12218 18163 12228 18316
rect 12334 18163 12344 18316
rect 12410 18163 12420 18316
rect 12456 18103 12676 18350
rect 12818 18163 12828 18316
rect 12894 18163 12904 18316
rect 13010 18163 13020 18316
rect 13086 18163 13096 18316
rect 13202 18163 13212 18316
rect 13278 18163 13288 18316
rect 13394 18163 13404 18316
rect 13470 18163 13480 18316
rect 13586 18163 13596 18316
rect 13662 18163 13672 18316
rect 13778 18163 13788 18316
rect 13854 18163 13864 18316
rect 13970 18163 13980 18316
rect 14046 18163 14056 18316
rect 14162 18163 14172 18316
rect 14238 18163 14248 18316
rect 14284 18103 14504 18350
rect 14646 18163 14656 18316
rect 14722 18163 14732 18316
rect 14838 18163 14848 18316
rect 14914 18163 14924 18316
rect 15030 18163 15040 18316
rect 15106 18163 15116 18316
rect 15222 18163 15232 18316
rect 15298 18163 15308 18316
rect 15414 18163 15424 18316
rect 15490 18163 15500 18316
rect 15606 18163 15616 18316
rect 15682 18163 15692 18316
rect 15798 18163 15808 18316
rect 15874 18163 15884 18316
rect 15990 18163 16000 18316
rect 16066 18163 16076 18316
rect 16112 18103 16332 18350
rect 16474 18163 16484 18316
rect 16550 18163 16560 18316
rect 16666 18163 16676 18316
rect 16742 18163 16752 18316
rect 16858 18163 16868 18316
rect 16934 18163 16944 18316
rect 17050 18163 17060 18316
rect 17126 18163 17136 18316
rect 17242 18163 17252 18316
rect 17318 18163 17328 18316
rect 17434 18163 17444 18316
rect 17510 18163 17520 18316
rect 17626 18163 17636 18316
rect 17702 18163 17712 18316
rect 17818 18163 17828 18316
rect 17894 18163 17904 18316
rect 17940 18103 18160 18350
rect 18302 18163 18312 18316
rect 18378 18163 18388 18316
rect 18494 18163 18504 18316
rect 18570 18163 18580 18316
rect 18686 18163 18696 18316
rect 18762 18163 18772 18316
rect 18878 18163 18888 18316
rect 18954 18163 18964 18316
rect 19070 18163 19080 18316
rect 19146 18163 19156 18316
rect 19262 18163 19272 18316
rect 19338 18163 19348 18316
rect 19454 18163 19464 18316
rect 19530 18163 19540 18316
rect 19646 18163 19656 18316
rect 19722 18163 19732 18316
rect 19768 18103 19988 18350
rect 20130 18163 20140 18316
rect 20206 18163 20216 18316
rect 20322 18163 20332 18316
rect 20398 18163 20408 18316
rect 20514 18163 20524 18316
rect 20590 18163 20600 18316
rect 20706 18163 20716 18316
rect 20782 18163 20792 18316
rect 20898 18163 20908 18316
rect 20974 18163 20984 18316
rect 21090 18163 21100 18316
rect 21166 18163 21176 18316
rect 21282 18163 21292 18316
rect 21358 18163 21368 18316
rect 21474 18163 21484 18316
rect 21550 18163 21560 18316
rect 21596 18103 21816 18350
rect 118 17950 128 18103
rect 194 17950 204 18103
rect 310 17950 320 18103
rect 386 17950 396 18103
rect 502 17950 512 18103
rect 578 17950 588 18103
rect 694 17950 704 18103
rect 770 17950 780 18103
rect 886 17950 896 18103
rect 962 17950 972 18103
rect 1078 17950 1088 18103
rect 1154 17950 1164 18103
rect 1270 17950 1280 18103
rect 1346 17950 1356 18103
rect 1462 17950 1472 18103
rect 1528 17950 1708 18103
rect 1946 17950 1956 18103
rect 2022 17950 2032 18103
rect 2138 17950 2148 18103
rect 2214 17950 2224 18103
rect 2330 17950 2340 18103
rect 2406 17950 2416 18103
rect 2522 17950 2532 18103
rect 2598 17950 2608 18103
rect 2714 17950 2724 18103
rect 2790 17950 2800 18103
rect 2906 17950 2916 18103
rect 2982 17950 2992 18103
rect 3098 17950 3108 18103
rect 3174 17950 3184 18103
rect 3290 17950 3300 18103
rect 3356 17950 3536 18103
rect 3774 17950 3784 18103
rect 3850 17950 3860 18103
rect 3966 17950 3976 18103
rect 4042 17950 4052 18103
rect 4158 17950 4168 18103
rect 4234 17950 4244 18103
rect 4350 17950 4360 18103
rect 4426 17950 4436 18103
rect 4542 17950 4552 18103
rect 4618 17950 4628 18103
rect 4734 17950 4744 18103
rect 4810 17950 4820 18103
rect 4926 17950 4936 18103
rect 5002 17950 5012 18103
rect 5118 17950 5128 18103
rect 5184 17950 5364 18103
rect 5602 17950 5612 18103
rect 5678 17950 5688 18103
rect 5794 17950 5804 18103
rect 5870 17950 5880 18103
rect 5986 17950 5996 18103
rect 6062 17950 6072 18103
rect 6178 17950 6188 18103
rect 6254 17950 6264 18103
rect 6370 17950 6380 18103
rect 6446 17950 6456 18103
rect 6562 17950 6572 18103
rect 6638 17950 6648 18103
rect 6754 17950 6764 18103
rect 6830 17950 6840 18103
rect 6946 17950 6956 18103
rect 7012 17950 7192 18103
rect 7430 17950 7440 18103
rect 7506 17950 7516 18103
rect 7622 17950 7632 18103
rect 7698 17950 7708 18103
rect 7814 17950 7824 18103
rect 7890 17950 7900 18103
rect 8006 17950 8016 18103
rect 8082 17950 8092 18103
rect 8198 17950 8208 18103
rect 8274 17950 8284 18103
rect 8390 17950 8400 18103
rect 8466 17950 8476 18103
rect 8582 17950 8592 18103
rect 8658 17950 8668 18103
rect 8774 17950 8784 18103
rect 8840 17950 9020 18103
rect 9258 17950 9268 18103
rect 9334 17950 9344 18103
rect 9450 17950 9460 18103
rect 9526 17950 9536 18103
rect 9642 17950 9652 18103
rect 9718 17950 9728 18103
rect 9834 17950 9844 18103
rect 9910 17950 9920 18103
rect 10026 17950 10036 18103
rect 10102 17950 10112 18103
rect 10218 17950 10228 18103
rect 10294 17950 10304 18103
rect 10410 17950 10420 18103
rect 10486 17950 10496 18103
rect 10602 17950 10612 18103
rect 10668 17950 10848 18103
rect 11086 17950 11096 18103
rect 11162 17950 11172 18103
rect 11278 17950 11288 18103
rect 11354 17950 11364 18103
rect 11470 17950 11480 18103
rect 11546 17950 11556 18103
rect 11662 17950 11672 18103
rect 11738 17950 11748 18103
rect 11854 17950 11864 18103
rect 11930 17950 11940 18103
rect 12046 17950 12056 18103
rect 12122 17950 12132 18103
rect 12238 17950 12248 18103
rect 12314 17950 12324 18103
rect 12430 17950 12440 18103
rect 12496 17950 12676 18103
rect 12914 17950 12924 18103
rect 12990 17950 13000 18103
rect 13106 17950 13116 18103
rect 13182 17950 13192 18103
rect 13298 17950 13308 18103
rect 13374 17950 13384 18103
rect 13490 17950 13500 18103
rect 13566 17950 13576 18103
rect 13682 17950 13692 18103
rect 13758 17950 13768 18103
rect 13874 17950 13884 18103
rect 13950 17950 13960 18103
rect 14066 17950 14076 18103
rect 14142 17950 14152 18103
rect 14258 17950 14268 18103
rect 14324 17950 14504 18103
rect 14742 17950 14752 18103
rect 14818 17950 14828 18103
rect 14934 17950 14944 18103
rect 15010 17950 15020 18103
rect 15126 17950 15136 18103
rect 15202 17950 15212 18103
rect 15318 17950 15328 18103
rect 15394 17950 15404 18103
rect 15510 17950 15520 18103
rect 15586 17950 15596 18103
rect 15702 17950 15712 18103
rect 15778 17950 15788 18103
rect 15894 17950 15904 18103
rect 15970 17950 15980 18103
rect 16086 17950 16096 18103
rect 16152 17950 16332 18103
rect 16570 17950 16580 18103
rect 16646 17950 16656 18103
rect 16762 17950 16772 18103
rect 16838 17950 16848 18103
rect 16954 17950 16964 18103
rect 17030 17950 17040 18103
rect 17146 17950 17156 18103
rect 17222 17950 17232 18103
rect 17338 17950 17348 18103
rect 17414 17950 17424 18103
rect 17530 17950 17540 18103
rect 17606 17950 17616 18103
rect 17722 17950 17732 18103
rect 17798 17950 17808 18103
rect 17914 17950 17924 18103
rect 17980 17950 18160 18103
rect 18398 17950 18408 18103
rect 18474 17950 18484 18103
rect 18590 17950 18600 18103
rect 18666 17950 18676 18103
rect 18782 17950 18792 18103
rect 18858 17950 18868 18103
rect 18974 17950 18984 18103
rect 19050 17950 19060 18103
rect 19166 17950 19176 18103
rect 19242 17950 19252 18103
rect 19358 17950 19368 18103
rect 19434 17950 19444 18103
rect 19550 17950 19560 18103
rect 19626 17950 19636 18103
rect 19742 17950 19752 18103
rect 19808 17950 19988 18103
rect 20226 17950 20236 18103
rect 20302 17950 20312 18103
rect 20418 17950 20428 18103
rect 20494 17950 20504 18103
rect 20610 17950 20620 18103
rect 20686 17950 20696 18103
rect 20802 17950 20812 18103
rect 20878 17950 20888 18103
rect 20994 17950 21004 18103
rect 21070 17950 21080 18103
rect 21186 17950 21196 18103
rect 21262 17950 21272 18103
rect 21378 17950 21388 18103
rect 21454 17950 21464 18103
rect 21570 17950 21580 18103
rect 21636 17950 21816 18103
rect 0 17853 1490 17912
rect 1828 17853 3318 17912
rect 3656 17853 5146 17912
rect 5484 17853 6974 17912
rect 7312 17853 8802 17912
rect 9140 17853 10630 17912
rect 10968 17853 12458 17912
rect 12796 17853 14286 17912
rect 14624 17853 16114 17912
rect 16452 17853 17942 17912
rect 18280 17853 19770 17912
rect 20108 17853 21598 17912
rect 0 17674 1490 17733
rect 1828 17674 3318 17733
rect 3656 17674 5146 17733
rect 5484 17674 6974 17733
rect 7312 17674 8802 17733
rect 9140 17674 10630 17733
rect 10968 17674 12458 17733
rect 12796 17674 14286 17733
rect 14624 17674 16114 17733
rect 16452 17674 17942 17733
rect 18280 17674 19770 17733
rect 20108 17674 21598 17733
rect 22 17449 32 17602
rect 98 17449 108 17602
rect 214 17449 224 17602
rect 290 17449 300 17602
rect 406 17449 416 17602
rect 482 17449 492 17602
rect 598 17449 608 17602
rect 674 17449 684 17602
rect 790 17449 800 17602
rect 866 17449 876 17602
rect 982 17449 992 17602
rect 1058 17449 1068 17602
rect 1174 17449 1184 17602
rect 1250 17449 1260 17602
rect 1366 17449 1376 17602
rect 1442 17449 1452 17602
rect 1488 17389 1708 17636
rect 1850 17449 1860 17602
rect 1926 17449 1936 17602
rect 2042 17449 2052 17602
rect 2118 17449 2128 17602
rect 2234 17449 2244 17602
rect 2310 17449 2320 17602
rect 2426 17449 2436 17602
rect 2502 17449 2512 17602
rect 2618 17449 2628 17602
rect 2694 17449 2704 17602
rect 2810 17449 2820 17602
rect 2886 17449 2896 17602
rect 3002 17449 3012 17602
rect 3078 17449 3088 17602
rect 3194 17449 3204 17602
rect 3270 17449 3280 17602
rect 3316 17389 3536 17636
rect 3678 17449 3688 17602
rect 3754 17449 3764 17602
rect 3870 17449 3880 17602
rect 3946 17449 3956 17602
rect 4062 17449 4072 17602
rect 4138 17449 4148 17602
rect 4254 17449 4264 17602
rect 4330 17449 4340 17602
rect 4446 17449 4456 17602
rect 4522 17449 4532 17602
rect 4638 17449 4648 17602
rect 4714 17449 4724 17602
rect 4830 17449 4840 17602
rect 4906 17449 4916 17602
rect 5022 17449 5032 17602
rect 5098 17449 5108 17602
rect 5144 17389 5364 17636
rect 5506 17449 5516 17602
rect 5582 17449 5592 17602
rect 5698 17449 5708 17602
rect 5774 17449 5784 17602
rect 5890 17449 5900 17602
rect 5966 17449 5976 17602
rect 6082 17449 6092 17602
rect 6158 17449 6168 17602
rect 6274 17449 6284 17602
rect 6350 17449 6360 17602
rect 6466 17449 6476 17602
rect 6542 17449 6552 17602
rect 6658 17449 6668 17602
rect 6734 17449 6744 17602
rect 6850 17449 6860 17602
rect 6926 17449 6936 17602
rect 6972 17389 7192 17636
rect 7334 17449 7344 17602
rect 7410 17449 7420 17602
rect 7526 17449 7536 17602
rect 7602 17449 7612 17602
rect 7718 17449 7728 17602
rect 7794 17449 7804 17602
rect 7910 17449 7920 17602
rect 7986 17449 7996 17602
rect 8102 17449 8112 17602
rect 8178 17449 8188 17602
rect 8294 17449 8304 17602
rect 8370 17449 8380 17602
rect 8486 17449 8496 17602
rect 8562 17449 8572 17602
rect 8678 17449 8688 17602
rect 8754 17449 8764 17602
rect 8800 17389 9020 17636
rect 9162 17449 9172 17602
rect 9238 17449 9248 17602
rect 9354 17449 9364 17602
rect 9430 17449 9440 17602
rect 9546 17449 9556 17602
rect 9622 17449 9632 17602
rect 9738 17449 9748 17602
rect 9814 17449 9824 17602
rect 9930 17449 9940 17602
rect 10006 17449 10016 17602
rect 10122 17449 10132 17602
rect 10198 17449 10208 17602
rect 10314 17449 10324 17602
rect 10390 17449 10400 17602
rect 10506 17449 10516 17602
rect 10582 17449 10592 17602
rect 10628 17389 10848 17636
rect 10990 17449 11000 17602
rect 11066 17449 11076 17602
rect 11182 17449 11192 17602
rect 11258 17449 11268 17602
rect 11374 17449 11384 17602
rect 11450 17449 11460 17602
rect 11566 17449 11576 17602
rect 11642 17449 11652 17602
rect 11758 17449 11768 17602
rect 11834 17449 11844 17602
rect 11950 17449 11960 17602
rect 12026 17449 12036 17602
rect 12142 17449 12152 17602
rect 12218 17449 12228 17602
rect 12334 17449 12344 17602
rect 12410 17449 12420 17602
rect 12456 17389 12676 17636
rect 12818 17449 12828 17602
rect 12894 17449 12904 17602
rect 13010 17449 13020 17602
rect 13086 17449 13096 17602
rect 13202 17449 13212 17602
rect 13278 17449 13288 17602
rect 13394 17449 13404 17602
rect 13470 17449 13480 17602
rect 13586 17449 13596 17602
rect 13662 17449 13672 17602
rect 13778 17449 13788 17602
rect 13854 17449 13864 17602
rect 13970 17449 13980 17602
rect 14046 17449 14056 17602
rect 14162 17449 14172 17602
rect 14238 17449 14248 17602
rect 14284 17389 14504 17636
rect 14646 17449 14656 17602
rect 14722 17449 14732 17602
rect 14838 17449 14848 17602
rect 14914 17449 14924 17602
rect 15030 17449 15040 17602
rect 15106 17449 15116 17602
rect 15222 17449 15232 17602
rect 15298 17449 15308 17602
rect 15414 17449 15424 17602
rect 15490 17449 15500 17602
rect 15606 17449 15616 17602
rect 15682 17449 15692 17602
rect 15798 17449 15808 17602
rect 15874 17449 15884 17602
rect 15990 17449 16000 17602
rect 16066 17449 16076 17602
rect 16112 17389 16332 17636
rect 16474 17449 16484 17602
rect 16550 17449 16560 17602
rect 16666 17449 16676 17602
rect 16742 17449 16752 17602
rect 16858 17449 16868 17602
rect 16934 17449 16944 17602
rect 17050 17449 17060 17602
rect 17126 17449 17136 17602
rect 17242 17449 17252 17602
rect 17318 17449 17328 17602
rect 17434 17449 17444 17602
rect 17510 17449 17520 17602
rect 17626 17449 17636 17602
rect 17702 17449 17712 17602
rect 17818 17449 17828 17602
rect 17894 17449 17904 17602
rect 17940 17389 18160 17636
rect 18302 17449 18312 17602
rect 18378 17449 18388 17602
rect 18494 17449 18504 17602
rect 18570 17449 18580 17602
rect 18686 17449 18696 17602
rect 18762 17449 18772 17602
rect 18878 17449 18888 17602
rect 18954 17449 18964 17602
rect 19070 17449 19080 17602
rect 19146 17449 19156 17602
rect 19262 17449 19272 17602
rect 19338 17449 19348 17602
rect 19454 17449 19464 17602
rect 19530 17449 19540 17602
rect 19646 17449 19656 17602
rect 19722 17449 19732 17602
rect 19768 17389 19988 17636
rect 20130 17449 20140 17602
rect 20206 17449 20216 17602
rect 20322 17449 20332 17602
rect 20398 17449 20408 17602
rect 20514 17449 20524 17602
rect 20590 17449 20600 17602
rect 20706 17449 20716 17602
rect 20782 17449 20792 17602
rect 20898 17449 20908 17602
rect 20974 17449 20984 17602
rect 21090 17449 21100 17602
rect 21166 17449 21176 17602
rect 21282 17449 21292 17602
rect 21358 17449 21368 17602
rect 21474 17449 21484 17602
rect 21550 17449 21560 17602
rect 21596 17389 21816 17636
rect 118 17236 128 17389
rect 194 17236 204 17389
rect 310 17236 320 17389
rect 386 17236 396 17389
rect 502 17236 512 17389
rect 578 17236 588 17389
rect 694 17236 704 17389
rect 770 17236 780 17389
rect 886 17236 896 17389
rect 962 17236 972 17389
rect 1078 17236 1088 17389
rect 1154 17236 1164 17389
rect 1270 17236 1280 17389
rect 1346 17236 1356 17389
rect 1462 17236 1472 17389
rect 1528 17236 1708 17389
rect 1946 17236 1956 17389
rect 2022 17236 2032 17389
rect 2138 17236 2148 17389
rect 2214 17236 2224 17389
rect 2330 17236 2340 17389
rect 2406 17236 2416 17389
rect 2522 17236 2532 17389
rect 2598 17236 2608 17389
rect 2714 17236 2724 17389
rect 2790 17236 2800 17389
rect 2906 17236 2916 17389
rect 2982 17236 2992 17389
rect 3098 17236 3108 17389
rect 3174 17236 3184 17389
rect 3290 17236 3300 17389
rect 3356 17236 3536 17389
rect 3774 17236 3784 17389
rect 3850 17236 3860 17389
rect 3966 17236 3976 17389
rect 4042 17236 4052 17389
rect 4158 17236 4168 17389
rect 4234 17236 4244 17389
rect 4350 17236 4360 17389
rect 4426 17236 4436 17389
rect 4542 17236 4552 17389
rect 4618 17236 4628 17389
rect 4734 17236 4744 17389
rect 4810 17236 4820 17389
rect 4926 17236 4936 17389
rect 5002 17236 5012 17389
rect 5118 17236 5128 17389
rect 5184 17236 5364 17389
rect 5602 17236 5612 17389
rect 5678 17236 5688 17389
rect 5794 17236 5804 17389
rect 5870 17236 5880 17389
rect 5986 17236 5996 17389
rect 6062 17236 6072 17389
rect 6178 17236 6188 17389
rect 6254 17236 6264 17389
rect 6370 17236 6380 17389
rect 6446 17236 6456 17389
rect 6562 17236 6572 17389
rect 6638 17236 6648 17389
rect 6754 17236 6764 17389
rect 6830 17236 6840 17389
rect 6946 17236 6956 17389
rect 7012 17236 7192 17389
rect 7430 17236 7440 17389
rect 7506 17236 7516 17389
rect 7622 17236 7632 17389
rect 7698 17236 7708 17389
rect 7814 17236 7824 17389
rect 7890 17236 7900 17389
rect 8006 17236 8016 17389
rect 8082 17236 8092 17389
rect 8198 17236 8208 17389
rect 8274 17236 8284 17389
rect 8390 17236 8400 17389
rect 8466 17236 8476 17389
rect 8582 17236 8592 17389
rect 8658 17236 8668 17389
rect 8774 17236 8784 17389
rect 8840 17236 9020 17389
rect 9258 17236 9268 17389
rect 9334 17236 9344 17389
rect 9450 17236 9460 17389
rect 9526 17236 9536 17389
rect 9642 17236 9652 17389
rect 9718 17236 9728 17389
rect 9834 17236 9844 17389
rect 9910 17236 9920 17389
rect 10026 17236 10036 17389
rect 10102 17236 10112 17389
rect 10218 17236 10228 17389
rect 10294 17236 10304 17389
rect 10410 17236 10420 17389
rect 10486 17236 10496 17389
rect 10602 17236 10612 17389
rect 10668 17236 10848 17389
rect 11086 17236 11096 17389
rect 11162 17236 11172 17389
rect 11278 17236 11288 17389
rect 11354 17236 11364 17389
rect 11470 17236 11480 17389
rect 11546 17236 11556 17389
rect 11662 17236 11672 17389
rect 11738 17236 11748 17389
rect 11854 17236 11864 17389
rect 11930 17236 11940 17389
rect 12046 17236 12056 17389
rect 12122 17236 12132 17389
rect 12238 17236 12248 17389
rect 12314 17236 12324 17389
rect 12430 17236 12440 17389
rect 12496 17236 12676 17389
rect 12914 17236 12924 17389
rect 12990 17236 13000 17389
rect 13106 17236 13116 17389
rect 13182 17236 13192 17389
rect 13298 17236 13308 17389
rect 13374 17236 13384 17389
rect 13490 17236 13500 17389
rect 13566 17236 13576 17389
rect 13682 17236 13692 17389
rect 13758 17236 13768 17389
rect 13874 17236 13884 17389
rect 13950 17236 13960 17389
rect 14066 17236 14076 17389
rect 14142 17236 14152 17389
rect 14258 17236 14268 17389
rect 14324 17236 14504 17389
rect 14742 17236 14752 17389
rect 14818 17236 14828 17389
rect 14934 17236 14944 17389
rect 15010 17236 15020 17389
rect 15126 17236 15136 17389
rect 15202 17236 15212 17389
rect 15318 17236 15328 17389
rect 15394 17236 15404 17389
rect 15510 17236 15520 17389
rect 15586 17236 15596 17389
rect 15702 17236 15712 17389
rect 15778 17236 15788 17389
rect 15894 17236 15904 17389
rect 15970 17236 15980 17389
rect 16086 17236 16096 17389
rect 16152 17236 16332 17389
rect 16570 17236 16580 17389
rect 16646 17236 16656 17389
rect 16762 17236 16772 17389
rect 16838 17236 16848 17389
rect 16954 17236 16964 17389
rect 17030 17236 17040 17389
rect 17146 17236 17156 17389
rect 17222 17236 17232 17389
rect 17338 17236 17348 17389
rect 17414 17236 17424 17389
rect 17530 17236 17540 17389
rect 17606 17236 17616 17389
rect 17722 17236 17732 17389
rect 17798 17236 17808 17389
rect 17914 17236 17924 17389
rect 17980 17236 18160 17389
rect 18398 17236 18408 17389
rect 18474 17236 18484 17389
rect 18590 17236 18600 17389
rect 18666 17236 18676 17389
rect 18782 17236 18792 17389
rect 18858 17236 18868 17389
rect 18974 17236 18984 17389
rect 19050 17236 19060 17389
rect 19166 17236 19176 17389
rect 19242 17236 19252 17389
rect 19358 17236 19368 17389
rect 19434 17236 19444 17389
rect 19550 17236 19560 17389
rect 19626 17236 19636 17389
rect 19742 17236 19752 17389
rect 19808 17236 19988 17389
rect 20226 17236 20236 17389
rect 20302 17236 20312 17389
rect 20418 17236 20428 17389
rect 20494 17236 20504 17389
rect 20610 17236 20620 17389
rect 20686 17236 20696 17389
rect 20802 17236 20812 17389
rect 20878 17236 20888 17389
rect 20994 17236 21004 17389
rect 21070 17236 21080 17389
rect 21186 17236 21196 17389
rect 21262 17236 21272 17389
rect 21378 17236 21388 17389
rect 21454 17236 21464 17389
rect 21570 17236 21580 17389
rect 21636 17236 21816 17389
rect 0 17139 1490 17198
rect 1828 17139 3318 17198
rect 3656 17139 5146 17198
rect 5484 17139 6974 17198
rect 7312 17139 8802 17198
rect 9140 17139 10630 17198
rect 10968 17139 12458 17198
rect 12796 17139 14286 17198
rect 14624 17139 16114 17198
rect 16452 17139 17942 17198
rect 18280 17139 19770 17198
rect 20108 17139 21598 17198
rect 0 16960 1490 17019
rect 1828 16960 3318 17019
rect 3656 16960 5146 17019
rect 5484 16960 6974 17019
rect 7312 16960 8802 17019
rect 9140 16960 10630 17019
rect 10968 16960 12458 17019
rect 12796 16960 14286 17019
rect 14624 16960 16114 17019
rect 16452 16960 17942 17019
rect 18280 16960 19770 17019
rect 20108 16960 21598 17019
rect 22 16735 32 16888
rect 98 16735 108 16888
rect 214 16735 224 16888
rect 290 16735 300 16888
rect 406 16735 416 16888
rect 482 16735 492 16888
rect 598 16735 608 16888
rect 674 16735 684 16888
rect 790 16735 800 16888
rect 866 16735 876 16888
rect 982 16735 992 16888
rect 1058 16735 1068 16888
rect 1174 16735 1184 16888
rect 1250 16735 1260 16888
rect 1366 16735 1376 16888
rect 1442 16735 1452 16888
rect 1488 16675 1708 16922
rect 1850 16735 1860 16888
rect 1926 16735 1936 16888
rect 2042 16735 2052 16888
rect 2118 16735 2128 16888
rect 2234 16735 2244 16888
rect 2310 16735 2320 16888
rect 2426 16735 2436 16888
rect 2502 16735 2512 16888
rect 2618 16735 2628 16888
rect 2694 16735 2704 16888
rect 2810 16735 2820 16888
rect 2886 16735 2896 16888
rect 3002 16735 3012 16888
rect 3078 16735 3088 16888
rect 3194 16735 3204 16888
rect 3270 16735 3280 16888
rect 3316 16675 3536 16922
rect 3678 16735 3688 16888
rect 3754 16735 3764 16888
rect 3870 16735 3880 16888
rect 3946 16735 3956 16888
rect 4062 16735 4072 16888
rect 4138 16735 4148 16888
rect 4254 16735 4264 16888
rect 4330 16735 4340 16888
rect 4446 16735 4456 16888
rect 4522 16735 4532 16888
rect 4638 16735 4648 16888
rect 4714 16735 4724 16888
rect 4830 16735 4840 16888
rect 4906 16735 4916 16888
rect 5022 16735 5032 16888
rect 5098 16735 5108 16888
rect 5144 16675 5364 16922
rect 5506 16735 5516 16888
rect 5582 16735 5592 16888
rect 5698 16735 5708 16888
rect 5774 16735 5784 16888
rect 5890 16735 5900 16888
rect 5966 16735 5976 16888
rect 6082 16735 6092 16888
rect 6158 16735 6168 16888
rect 6274 16735 6284 16888
rect 6350 16735 6360 16888
rect 6466 16735 6476 16888
rect 6542 16735 6552 16888
rect 6658 16735 6668 16888
rect 6734 16735 6744 16888
rect 6850 16735 6860 16888
rect 6926 16735 6936 16888
rect 6972 16675 7192 16922
rect 7334 16735 7344 16888
rect 7410 16735 7420 16888
rect 7526 16735 7536 16888
rect 7602 16735 7612 16888
rect 7718 16735 7728 16888
rect 7794 16735 7804 16888
rect 7910 16735 7920 16888
rect 7986 16735 7996 16888
rect 8102 16735 8112 16888
rect 8178 16735 8188 16888
rect 8294 16735 8304 16888
rect 8370 16735 8380 16888
rect 8486 16735 8496 16888
rect 8562 16735 8572 16888
rect 8678 16735 8688 16888
rect 8754 16735 8764 16888
rect 8800 16675 9020 16922
rect 9162 16735 9172 16888
rect 9238 16735 9248 16888
rect 9354 16735 9364 16888
rect 9430 16735 9440 16888
rect 9546 16735 9556 16888
rect 9622 16735 9632 16888
rect 9738 16735 9748 16888
rect 9814 16735 9824 16888
rect 9930 16735 9940 16888
rect 10006 16735 10016 16888
rect 10122 16735 10132 16888
rect 10198 16735 10208 16888
rect 10314 16735 10324 16888
rect 10390 16735 10400 16888
rect 10506 16735 10516 16888
rect 10582 16735 10592 16888
rect 10628 16675 10848 16922
rect 10990 16735 11000 16888
rect 11066 16735 11076 16888
rect 11182 16735 11192 16888
rect 11258 16735 11268 16888
rect 11374 16735 11384 16888
rect 11450 16735 11460 16888
rect 11566 16735 11576 16888
rect 11642 16735 11652 16888
rect 11758 16735 11768 16888
rect 11834 16735 11844 16888
rect 11950 16735 11960 16888
rect 12026 16735 12036 16888
rect 12142 16735 12152 16888
rect 12218 16735 12228 16888
rect 12334 16735 12344 16888
rect 12410 16735 12420 16888
rect 12456 16675 12676 16922
rect 12818 16735 12828 16888
rect 12894 16735 12904 16888
rect 13010 16735 13020 16888
rect 13086 16735 13096 16888
rect 13202 16735 13212 16888
rect 13278 16735 13288 16888
rect 13394 16735 13404 16888
rect 13470 16735 13480 16888
rect 13586 16735 13596 16888
rect 13662 16735 13672 16888
rect 13778 16735 13788 16888
rect 13854 16735 13864 16888
rect 13970 16735 13980 16888
rect 14046 16735 14056 16888
rect 14162 16735 14172 16888
rect 14238 16735 14248 16888
rect 14284 16675 14504 16922
rect 14646 16735 14656 16888
rect 14722 16735 14732 16888
rect 14838 16735 14848 16888
rect 14914 16735 14924 16888
rect 15030 16735 15040 16888
rect 15106 16735 15116 16888
rect 15222 16735 15232 16888
rect 15298 16735 15308 16888
rect 15414 16735 15424 16888
rect 15490 16735 15500 16888
rect 15606 16735 15616 16888
rect 15682 16735 15692 16888
rect 15798 16735 15808 16888
rect 15874 16735 15884 16888
rect 15990 16735 16000 16888
rect 16066 16735 16076 16888
rect 16112 16675 16332 16922
rect 16474 16735 16484 16888
rect 16550 16735 16560 16888
rect 16666 16735 16676 16888
rect 16742 16735 16752 16888
rect 16858 16735 16868 16888
rect 16934 16735 16944 16888
rect 17050 16735 17060 16888
rect 17126 16735 17136 16888
rect 17242 16735 17252 16888
rect 17318 16735 17328 16888
rect 17434 16735 17444 16888
rect 17510 16735 17520 16888
rect 17626 16735 17636 16888
rect 17702 16735 17712 16888
rect 17818 16735 17828 16888
rect 17894 16735 17904 16888
rect 17940 16675 18160 16922
rect 18302 16735 18312 16888
rect 18378 16735 18388 16888
rect 18494 16735 18504 16888
rect 18570 16735 18580 16888
rect 18686 16735 18696 16888
rect 18762 16735 18772 16888
rect 18878 16735 18888 16888
rect 18954 16735 18964 16888
rect 19070 16735 19080 16888
rect 19146 16735 19156 16888
rect 19262 16735 19272 16888
rect 19338 16735 19348 16888
rect 19454 16735 19464 16888
rect 19530 16735 19540 16888
rect 19646 16735 19656 16888
rect 19722 16735 19732 16888
rect 19768 16675 19988 16922
rect 20130 16735 20140 16888
rect 20206 16735 20216 16888
rect 20322 16735 20332 16888
rect 20398 16735 20408 16888
rect 20514 16735 20524 16888
rect 20590 16735 20600 16888
rect 20706 16735 20716 16888
rect 20782 16735 20792 16888
rect 20898 16735 20908 16888
rect 20974 16735 20984 16888
rect 21090 16735 21100 16888
rect 21166 16735 21176 16888
rect 21282 16735 21292 16888
rect 21358 16735 21368 16888
rect 21474 16735 21484 16888
rect 21550 16735 21560 16888
rect 21596 16675 21816 16922
rect 118 16522 128 16675
rect 194 16522 204 16675
rect 310 16522 320 16675
rect 386 16522 396 16675
rect 502 16522 512 16675
rect 578 16522 588 16675
rect 694 16522 704 16675
rect 770 16522 780 16675
rect 886 16522 896 16675
rect 962 16522 972 16675
rect 1078 16522 1088 16675
rect 1154 16522 1164 16675
rect 1270 16522 1280 16675
rect 1346 16522 1356 16675
rect 1462 16522 1472 16675
rect 1528 16522 1708 16675
rect 1946 16522 1956 16675
rect 2022 16522 2032 16675
rect 2138 16522 2148 16675
rect 2214 16522 2224 16675
rect 2330 16522 2340 16675
rect 2406 16522 2416 16675
rect 2522 16522 2532 16675
rect 2598 16522 2608 16675
rect 2714 16522 2724 16675
rect 2790 16522 2800 16675
rect 2906 16522 2916 16675
rect 2982 16522 2992 16675
rect 3098 16522 3108 16675
rect 3174 16522 3184 16675
rect 3290 16522 3300 16675
rect 3356 16522 3536 16675
rect 3774 16522 3784 16675
rect 3850 16522 3860 16675
rect 3966 16522 3976 16675
rect 4042 16522 4052 16675
rect 4158 16522 4168 16675
rect 4234 16522 4244 16675
rect 4350 16522 4360 16675
rect 4426 16522 4436 16675
rect 4542 16522 4552 16675
rect 4618 16522 4628 16675
rect 4734 16522 4744 16675
rect 4810 16522 4820 16675
rect 4926 16522 4936 16675
rect 5002 16522 5012 16675
rect 5118 16522 5128 16675
rect 5184 16522 5364 16675
rect 5602 16522 5612 16675
rect 5678 16522 5688 16675
rect 5794 16522 5804 16675
rect 5870 16522 5880 16675
rect 5986 16522 5996 16675
rect 6062 16522 6072 16675
rect 6178 16522 6188 16675
rect 6254 16522 6264 16675
rect 6370 16522 6380 16675
rect 6446 16522 6456 16675
rect 6562 16522 6572 16675
rect 6638 16522 6648 16675
rect 6754 16522 6764 16675
rect 6830 16522 6840 16675
rect 6946 16522 6956 16675
rect 7012 16522 7192 16675
rect 7430 16522 7440 16675
rect 7506 16522 7516 16675
rect 7622 16522 7632 16675
rect 7698 16522 7708 16675
rect 7814 16522 7824 16675
rect 7890 16522 7900 16675
rect 8006 16522 8016 16675
rect 8082 16522 8092 16675
rect 8198 16522 8208 16675
rect 8274 16522 8284 16675
rect 8390 16522 8400 16675
rect 8466 16522 8476 16675
rect 8582 16522 8592 16675
rect 8658 16522 8668 16675
rect 8774 16522 8784 16675
rect 8840 16522 9020 16675
rect 9258 16522 9268 16675
rect 9334 16522 9344 16675
rect 9450 16522 9460 16675
rect 9526 16522 9536 16675
rect 9642 16522 9652 16675
rect 9718 16522 9728 16675
rect 9834 16522 9844 16675
rect 9910 16522 9920 16675
rect 10026 16522 10036 16675
rect 10102 16522 10112 16675
rect 10218 16522 10228 16675
rect 10294 16522 10304 16675
rect 10410 16522 10420 16675
rect 10486 16522 10496 16675
rect 10602 16522 10612 16675
rect 10668 16522 10848 16675
rect 11086 16522 11096 16675
rect 11162 16522 11172 16675
rect 11278 16522 11288 16675
rect 11354 16522 11364 16675
rect 11470 16522 11480 16675
rect 11546 16522 11556 16675
rect 11662 16522 11672 16675
rect 11738 16522 11748 16675
rect 11854 16522 11864 16675
rect 11930 16522 11940 16675
rect 12046 16522 12056 16675
rect 12122 16522 12132 16675
rect 12238 16522 12248 16675
rect 12314 16522 12324 16675
rect 12430 16522 12440 16675
rect 12496 16522 12676 16675
rect 12914 16522 12924 16675
rect 12990 16522 13000 16675
rect 13106 16522 13116 16675
rect 13182 16522 13192 16675
rect 13298 16522 13308 16675
rect 13374 16522 13384 16675
rect 13490 16522 13500 16675
rect 13566 16522 13576 16675
rect 13682 16522 13692 16675
rect 13758 16522 13768 16675
rect 13874 16522 13884 16675
rect 13950 16522 13960 16675
rect 14066 16522 14076 16675
rect 14142 16522 14152 16675
rect 14258 16522 14268 16675
rect 14324 16522 14504 16675
rect 14742 16522 14752 16675
rect 14818 16522 14828 16675
rect 14934 16522 14944 16675
rect 15010 16522 15020 16675
rect 15126 16522 15136 16675
rect 15202 16522 15212 16675
rect 15318 16522 15328 16675
rect 15394 16522 15404 16675
rect 15510 16522 15520 16675
rect 15586 16522 15596 16675
rect 15702 16522 15712 16675
rect 15778 16522 15788 16675
rect 15894 16522 15904 16675
rect 15970 16522 15980 16675
rect 16086 16522 16096 16675
rect 16152 16522 16332 16675
rect 16570 16522 16580 16675
rect 16646 16522 16656 16675
rect 16762 16522 16772 16675
rect 16838 16522 16848 16675
rect 16954 16522 16964 16675
rect 17030 16522 17040 16675
rect 17146 16522 17156 16675
rect 17222 16522 17232 16675
rect 17338 16522 17348 16675
rect 17414 16522 17424 16675
rect 17530 16522 17540 16675
rect 17606 16522 17616 16675
rect 17722 16522 17732 16675
rect 17798 16522 17808 16675
rect 17914 16522 17924 16675
rect 17980 16522 18160 16675
rect 18398 16522 18408 16675
rect 18474 16522 18484 16675
rect 18590 16522 18600 16675
rect 18666 16522 18676 16675
rect 18782 16522 18792 16675
rect 18858 16522 18868 16675
rect 18974 16522 18984 16675
rect 19050 16522 19060 16675
rect 19166 16522 19176 16675
rect 19242 16522 19252 16675
rect 19358 16522 19368 16675
rect 19434 16522 19444 16675
rect 19550 16522 19560 16675
rect 19626 16522 19636 16675
rect 19742 16522 19752 16675
rect 19808 16522 19988 16675
rect 20226 16522 20236 16675
rect 20302 16522 20312 16675
rect 20418 16522 20428 16675
rect 20494 16522 20504 16675
rect 20610 16522 20620 16675
rect 20686 16522 20696 16675
rect 20802 16522 20812 16675
rect 20878 16522 20888 16675
rect 20994 16522 21004 16675
rect 21070 16522 21080 16675
rect 21186 16522 21196 16675
rect 21262 16522 21272 16675
rect 21378 16522 21388 16675
rect 21454 16522 21464 16675
rect 21570 16522 21580 16675
rect 21636 16522 21816 16675
rect 0 16425 1490 16484
rect 1828 16425 3318 16484
rect 3656 16425 5146 16484
rect 5484 16425 6974 16484
rect 7312 16425 8802 16484
rect 9140 16425 10630 16484
rect 10968 16425 12458 16484
rect 12796 16425 14286 16484
rect 14624 16425 16114 16484
rect 16452 16425 17942 16484
rect 18280 16425 19770 16484
rect 20108 16425 21598 16484
rect 0 16246 1490 16305
rect 1828 16246 3318 16305
rect 3656 16246 5146 16305
rect 5484 16246 6974 16305
rect 7312 16246 8802 16305
rect 9140 16246 10630 16305
rect 10968 16246 12458 16305
rect 12796 16246 14286 16305
rect 14624 16246 16114 16305
rect 16452 16246 17942 16305
rect 18280 16246 19770 16305
rect 20108 16246 21598 16305
rect 22 16021 32 16174
rect 98 16021 108 16174
rect 214 16021 224 16174
rect 290 16021 300 16174
rect 406 16021 416 16174
rect 482 16021 492 16174
rect 598 16021 608 16174
rect 674 16021 684 16174
rect 790 16021 800 16174
rect 866 16021 876 16174
rect 982 16021 992 16174
rect 1058 16021 1068 16174
rect 1174 16021 1184 16174
rect 1250 16021 1260 16174
rect 1366 16021 1376 16174
rect 1442 16021 1452 16174
rect 1488 15961 1708 16208
rect 1850 16021 1860 16174
rect 1926 16021 1936 16174
rect 2042 16021 2052 16174
rect 2118 16021 2128 16174
rect 2234 16021 2244 16174
rect 2310 16021 2320 16174
rect 2426 16021 2436 16174
rect 2502 16021 2512 16174
rect 2618 16021 2628 16174
rect 2694 16021 2704 16174
rect 2810 16021 2820 16174
rect 2886 16021 2896 16174
rect 3002 16021 3012 16174
rect 3078 16021 3088 16174
rect 3194 16021 3204 16174
rect 3270 16021 3280 16174
rect 3316 15961 3536 16208
rect 3678 16021 3688 16174
rect 3754 16021 3764 16174
rect 3870 16021 3880 16174
rect 3946 16021 3956 16174
rect 4062 16021 4072 16174
rect 4138 16021 4148 16174
rect 4254 16021 4264 16174
rect 4330 16021 4340 16174
rect 4446 16021 4456 16174
rect 4522 16021 4532 16174
rect 4638 16021 4648 16174
rect 4714 16021 4724 16174
rect 4830 16021 4840 16174
rect 4906 16021 4916 16174
rect 5022 16021 5032 16174
rect 5098 16021 5108 16174
rect 5144 15961 5364 16208
rect 5506 16021 5516 16174
rect 5582 16021 5592 16174
rect 5698 16021 5708 16174
rect 5774 16021 5784 16174
rect 5890 16021 5900 16174
rect 5966 16021 5976 16174
rect 6082 16021 6092 16174
rect 6158 16021 6168 16174
rect 6274 16021 6284 16174
rect 6350 16021 6360 16174
rect 6466 16021 6476 16174
rect 6542 16021 6552 16174
rect 6658 16021 6668 16174
rect 6734 16021 6744 16174
rect 6850 16021 6860 16174
rect 6926 16021 6936 16174
rect 6972 15961 7192 16208
rect 7334 16021 7344 16174
rect 7410 16021 7420 16174
rect 7526 16021 7536 16174
rect 7602 16021 7612 16174
rect 7718 16021 7728 16174
rect 7794 16021 7804 16174
rect 7910 16021 7920 16174
rect 7986 16021 7996 16174
rect 8102 16021 8112 16174
rect 8178 16021 8188 16174
rect 8294 16021 8304 16174
rect 8370 16021 8380 16174
rect 8486 16021 8496 16174
rect 8562 16021 8572 16174
rect 8678 16021 8688 16174
rect 8754 16021 8764 16174
rect 8800 15961 9020 16208
rect 9162 16021 9172 16174
rect 9238 16021 9248 16174
rect 9354 16021 9364 16174
rect 9430 16021 9440 16174
rect 9546 16021 9556 16174
rect 9622 16021 9632 16174
rect 9738 16021 9748 16174
rect 9814 16021 9824 16174
rect 9930 16021 9940 16174
rect 10006 16021 10016 16174
rect 10122 16021 10132 16174
rect 10198 16021 10208 16174
rect 10314 16021 10324 16174
rect 10390 16021 10400 16174
rect 10506 16021 10516 16174
rect 10582 16021 10592 16174
rect 10628 15961 10848 16208
rect 10990 16021 11000 16174
rect 11066 16021 11076 16174
rect 11182 16021 11192 16174
rect 11258 16021 11268 16174
rect 11374 16021 11384 16174
rect 11450 16021 11460 16174
rect 11566 16021 11576 16174
rect 11642 16021 11652 16174
rect 11758 16021 11768 16174
rect 11834 16021 11844 16174
rect 11950 16021 11960 16174
rect 12026 16021 12036 16174
rect 12142 16021 12152 16174
rect 12218 16021 12228 16174
rect 12334 16021 12344 16174
rect 12410 16021 12420 16174
rect 12456 15961 12676 16208
rect 12818 16021 12828 16174
rect 12894 16021 12904 16174
rect 13010 16021 13020 16174
rect 13086 16021 13096 16174
rect 13202 16021 13212 16174
rect 13278 16021 13288 16174
rect 13394 16021 13404 16174
rect 13470 16021 13480 16174
rect 13586 16021 13596 16174
rect 13662 16021 13672 16174
rect 13778 16021 13788 16174
rect 13854 16021 13864 16174
rect 13970 16021 13980 16174
rect 14046 16021 14056 16174
rect 14162 16021 14172 16174
rect 14238 16021 14248 16174
rect 14284 15961 14504 16208
rect 14646 16021 14656 16174
rect 14722 16021 14732 16174
rect 14838 16021 14848 16174
rect 14914 16021 14924 16174
rect 15030 16021 15040 16174
rect 15106 16021 15116 16174
rect 15222 16021 15232 16174
rect 15298 16021 15308 16174
rect 15414 16021 15424 16174
rect 15490 16021 15500 16174
rect 15606 16021 15616 16174
rect 15682 16021 15692 16174
rect 15798 16021 15808 16174
rect 15874 16021 15884 16174
rect 15990 16021 16000 16174
rect 16066 16021 16076 16174
rect 16112 15961 16332 16208
rect 16474 16021 16484 16174
rect 16550 16021 16560 16174
rect 16666 16021 16676 16174
rect 16742 16021 16752 16174
rect 16858 16021 16868 16174
rect 16934 16021 16944 16174
rect 17050 16021 17060 16174
rect 17126 16021 17136 16174
rect 17242 16021 17252 16174
rect 17318 16021 17328 16174
rect 17434 16021 17444 16174
rect 17510 16021 17520 16174
rect 17626 16021 17636 16174
rect 17702 16021 17712 16174
rect 17818 16021 17828 16174
rect 17894 16021 17904 16174
rect 17940 15961 18160 16208
rect 18302 16021 18312 16174
rect 18378 16021 18388 16174
rect 18494 16021 18504 16174
rect 18570 16021 18580 16174
rect 18686 16021 18696 16174
rect 18762 16021 18772 16174
rect 18878 16021 18888 16174
rect 18954 16021 18964 16174
rect 19070 16021 19080 16174
rect 19146 16021 19156 16174
rect 19262 16021 19272 16174
rect 19338 16021 19348 16174
rect 19454 16021 19464 16174
rect 19530 16021 19540 16174
rect 19646 16021 19656 16174
rect 19722 16021 19732 16174
rect 19768 15961 19988 16208
rect 20130 16021 20140 16174
rect 20206 16021 20216 16174
rect 20322 16021 20332 16174
rect 20398 16021 20408 16174
rect 20514 16021 20524 16174
rect 20590 16021 20600 16174
rect 20706 16021 20716 16174
rect 20782 16021 20792 16174
rect 20898 16021 20908 16174
rect 20974 16021 20984 16174
rect 21090 16021 21100 16174
rect 21166 16021 21176 16174
rect 21282 16021 21292 16174
rect 21358 16021 21368 16174
rect 21474 16021 21484 16174
rect 21550 16021 21560 16174
rect 21596 15961 21816 16208
rect 118 15808 128 15961
rect 194 15808 204 15961
rect 310 15808 320 15961
rect 386 15808 396 15961
rect 502 15808 512 15961
rect 578 15808 588 15961
rect 694 15808 704 15961
rect 770 15808 780 15961
rect 886 15808 896 15961
rect 962 15808 972 15961
rect 1078 15808 1088 15961
rect 1154 15808 1164 15961
rect 1270 15808 1280 15961
rect 1346 15808 1356 15961
rect 1462 15808 1472 15961
rect 1528 15808 1708 15961
rect 1946 15808 1956 15961
rect 2022 15808 2032 15961
rect 2138 15808 2148 15961
rect 2214 15808 2224 15961
rect 2330 15808 2340 15961
rect 2406 15808 2416 15961
rect 2522 15808 2532 15961
rect 2598 15808 2608 15961
rect 2714 15808 2724 15961
rect 2790 15808 2800 15961
rect 2906 15808 2916 15961
rect 2982 15808 2992 15961
rect 3098 15808 3108 15961
rect 3174 15808 3184 15961
rect 3290 15808 3300 15961
rect 3356 15808 3536 15961
rect 3774 15808 3784 15961
rect 3850 15808 3860 15961
rect 3966 15808 3976 15961
rect 4042 15808 4052 15961
rect 4158 15808 4168 15961
rect 4234 15808 4244 15961
rect 4350 15808 4360 15961
rect 4426 15808 4436 15961
rect 4542 15808 4552 15961
rect 4618 15808 4628 15961
rect 4734 15808 4744 15961
rect 4810 15808 4820 15961
rect 4926 15808 4936 15961
rect 5002 15808 5012 15961
rect 5118 15808 5128 15961
rect 5184 15808 5364 15961
rect 5602 15808 5612 15961
rect 5678 15808 5688 15961
rect 5794 15808 5804 15961
rect 5870 15808 5880 15961
rect 5986 15808 5996 15961
rect 6062 15808 6072 15961
rect 6178 15808 6188 15961
rect 6254 15808 6264 15961
rect 6370 15808 6380 15961
rect 6446 15808 6456 15961
rect 6562 15808 6572 15961
rect 6638 15808 6648 15961
rect 6754 15808 6764 15961
rect 6830 15808 6840 15961
rect 6946 15808 6956 15961
rect 7012 15808 7192 15961
rect 7430 15808 7440 15961
rect 7506 15808 7516 15961
rect 7622 15808 7632 15961
rect 7698 15808 7708 15961
rect 7814 15808 7824 15961
rect 7890 15808 7900 15961
rect 8006 15808 8016 15961
rect 8082 15808 8092 15961
rect 8198 15808 8208 15961
rect 8274 15808 8284 15961
rect 8390 15808 8400 15961
rect 8466 15808 8476 15961
rect 8582 15808 8592 15961
rect 8658 15808 8668 15961
rect 8774 15808 8784 15961
rect 8840 15808 9020 15961
rect 9258 15808 9268 15961
rect 9334 15808 9344 15961
rect 9450 15808 9460 15961
rect 9526 15808 9536 15961
rect 9642 15808 9652 15961
rect 9718 15808 9728 15961
rect 9834 15808 9844 15961
rect 9910 15808 9920 15961
rect 10026 15808 10036 15961
rect 10102 15808 10112 15961
rect 10218 15808 10228 15961
rect 10294 15808 10304 15961
rect 10410 15808 10420 15961
rect 10486 15808 10496 15961
rect 10602 15808 10612 15961
rect 10668 15808 10848 15961
rect 11086 15808 11096 15961
rect 11162 15808 11172 15961
rect 11278 15808 11288 15961
rect 11354 15808 11364 15961
rect 11470 15808 11480 15961
rect 11546 15808 11556 15961
rect 11662 15808 11672 15961
rect 11738 15808 11748 15961
rect 11854 15808 11864 15961
rect 11930 15808 11940 15961
rect 12046 15808 12056 15961
rect 12122 15808 12132 15961
rect 12238 15808 12248 15961
rect 12314 15808 12324 15961
rect 12430 15808 12440 15961
rect 12496 15808 12676 15961
rect 12914 15808 12924 15961
rect 12990 15808 13000 15961
rect 13106 15808 13116 15961
rect 13182 15808 13192 15961
rect 13298 15808 13308 15961
rect 13374 15808 13384 15961
rect 13490 15808 13500 15961
rect 13566 15808 13576 15961
rect 13682 15808 13692 15961
rect 13758 15808 13768 15961
rect 13874 15808 13884 15961
rect 13950 15808 13960 15961
rect 14066 15808 14076 15961
rect 14142 15808 14152 15961
rect 14258 15808 14268 15961
rect 14324 15808 14504 15961
rect 14742 15808 14752 15961
rect 14818 15808 14828 15961
rect 14934 15808 14944 15961
rect 15010 15808 15020 15961
rect 15126 15808 15136 15961
rect 15202 15808 15212 15961
rect 15318 15808 15328 15961
rect 15394 15808 15404 15961
rect 15510 15808 15520 15961
rect 15586 15808 15596 15961
rect 15702 15808 15712 15961
rect 15778 15808 15788 15961
rect 15894 15808 15904 15961
rect 15970 15808 15980 15961
rect 16086 15808 16096 15961
rect 16152 15808 16332 15961
rect 16570 15808 16580 15961
rect 16646 15808 16656 15961
rect 16762 15808 16772 15961
rect 16838 15808 16848 15961
rect 16954 15808 16964 15961
rect 17030 15808 17040 15961
rect 17146 15808 17156 15961
rect 17222 15808 17232 15961
rect 17338 15808 17348 15961
rect 17414 15808 17424 15961
rect 17530 15808 17540 15961
rect 17606 15808 17616 15961
rect 17722 15808 17732 15961
rect 17798 15808 17808 15961
rect 17914 15808 17924 15961
rect 17980 15808 18160 15961
rect 18398 15808 18408 15961
rect 18474 15808 18484 15961
rect 18590 15808 18600 15961
rect 18666 15808 18676 15961
rect 18782 15808 18792 15961
rect 18858 15808 18868 15961
rect 18974 15808 18984 15961
rect 19050 15808 19060 15961
rect 19166 15808 19176 15961
rect 19242 15808 19252 15961
rect 19358 15808 19368 15961
rect 19434 15808 19444 15961
rect 19550 15808 19560 15961
rect 19626 15808 19636 15961
rect 19742 15808 19752 15961
rect 19808 15808 19988 15961
rect 20226 15808 20236 15961
rect 20302 15808 20312 15961
rect 20418 15808 20428 15961
rect 20494 15808 20504 15961
rect 20610 15808 20620 15961
rect 20686 15808 20696 15961
rect 20802 15808 20812 15961
rect 20878 15808 20888 15961
rect 20994 15808 21004 15961
rect 21070 15808 21080 15961
rect 21186 15808 21196 15961
rect 21262 15808 21272 15961
rect 21378 15808 21388 15961
rect 21454 15808 21464 15961
rect 21570 15808 21580 15961
rect 21636 15808 21816 15961
rect 0 15711 1490 15770
rect 1828 15711 3318 15770
rect 3656 15711 5146 15770
rect 5484 15711 6974 15770
rect 7312 15711 8802 15770
rect 9140 15711 10630 15770
rect 10968 15711 12458 15770
rect 12796 15711 14286 15770
rect 14624 15711 16114 15770
rect 16452 15711 17942 15770
rect 18280 15711 19770 15770
rect 20108 15711 21598 15770
rect 0 15532 1490 15591
rect 1828 15532 3318 15591
rect 3656 15532 5146 15591
rect 5484 15532 6974 15591
rect 7312 15532 8802 15591
rect 9140 15532 10630 15591
rect 10968 15532 12458 15591
rect 12796 15532 14286 15591
rect 14624 15532 16114 15591
rect 16452 15532 17942 15591
rect 18280 15532 19770 15591
rect 20108 15532 21598 15591
rect 22 15307 32 15460
rect 98 15307 108 15460
rect 214 15307 224 15460
rect 290 15307 300 15460
rect 406 15307 416 15460
rect 482 15307 492 15460
rect 598 15307 608 15460
rect 674 15307 684 15460
rect 790 15307 800 15460
rect 866 15307 876 15460
rect 982 15307 992 15460
rect 1058 15307 1068 15460
rect 1174 15307 1184 15460
rect 1250 15307 1260 15460
rect 1366 15307 1376 15460
rect 1442 15307 1452 15460
rect 1488 15247 1708 15494
rect 1850 15307 1860 15460
rect 1926 15307 1936 15460
rect 2042 15307 2052 15460
rect 2118 15307 2128 15460
rect 2234 15307 2244 15460
rect 2310 15307 2320 15460
rect 2426 15307 2436 15460
rect 2502 15307 2512 15460
rect 2618 15307 2628 15460
rect 2694 15307 2704 15460
rect 2810 15307 2820 15460
rect 2886 15307 2896 15460
rect 3002 15307 3012 15460
rect 3078 15307 3088 15460
rect 3194 15307 3204 15460
rect 3270 15307 3280 15460
rect 3316 15247 3536 15494
rect 3678 15307 3688 15460
rect 3754 15307 3764 15460
rect 3870 15307 3880 15460
rect 3946 15307 3956 15460
rect 4062 15307 4072 15460
rect 4138 15307 4148 15460
rect 4254 15307 4264 15460
rect 4330 15307 4340 15460
rect 4446 15307 4456 15460
rect 4522 15307 4532 15460
rect 4638 15307 4648 15460
rect 4714 15307 4724 15460
rect 4830 15307 4840 15460
rect 4906 15307 4916 15460
rect 5022 15307 5032 15460
rect 5098 15307 5108 15460
rect 5144 15247 5364 15494
rect 5506 15307 5516 15460
rect 5582 15307 5592 15460
rect 5698 15307 5708 15460
rect 5774 15307 5784 15460
rect 5890 15307 5900 15460
rect 5966 15307 5976 15460
rect 6082 15307 6092 15460
rect 6158 15307 6168 15460
rect 6274 15307 6284 15460
rect 6350 15307 6360 15460
rect 6466 15307 6476 15460
rect 6542 15307 6552 15460
rect 6658 15307 6668 15460
rect 6734 15307 6744 15460
rect 6850 15307 6860 15460
rect 6926 15307 6936 15460
rect 6972 15247 7192 15494
rect 7334 15307 7344 15460
rect 7410 15307 7420 15460
rect 7526 15307 7536 15460
rect 7602 15307 7612 15460
rect 7718 15307 7728 15460
rect 7794 15307 7804 15460
rect 7910 15307 7920 15460
rect 7986 15307 7996 15460
rect 8102 15307 8112 15460
rect 8178 15307 8188 15460
rect 8294 15307 8304 15460
rect 8370 15307 8380 15460
rect 8486 15307 8496 15460
rect 8562 15307 8572 15460
rect 8678 15307 8688 15460
rect 8754 15307 8764 15460
rect 8800 15247 9020 15494
rect 9162 15307 9172 15460
rect 9238 15307 9248 15460
rect 9354 15307 9364 15460
rect 9430 15307 9440 15460
rect 9546 15307 9556 15460
rect 9622 15307 9632 15460
rect 9738 15307 9748 15460
rect 9814 15307 9824 15460
rect 9930 15307 9940 15460
rect 10006 15307 10016 15460
rect 10122 15307 10132 15460
rect 10198 15307 10208 15460
rect 10314 15307 10324 15460
rect 10390 15307 10400 15460
rect 10506 15307 10516 15460
rect 10582 15307 10592 15460
rect 10628 15247 10848 15494
rect 10990 15307 11000 15460
rect 11066 15307 11076 15460
rect 11182 15307 11192 15460
rect 11258 15307 11268 15460
rect 11374 15307 11384 15460
rect 11450 15307 11460 15460
rect 11566 15307 11576 15460
rect 11642 15307 11652 15460
rect 11758 15307 11768 15460
rect 11834 15307 11844 15460
rect 11950 15307 11960 15460
rect 12026 15307 12036 15460
rect 12142 15307 12152 15460
rect 12218 15307 12228 15460
rect 12334 15307 12344 15460
rect 12410 15307 12420 15460
rect 12456 15247 12676 15494
rect 12818 15307 12828 15460
rect 12894 15307 12904 15460
rect 13010 15307 13020 15460
rect 13086 15307 13096 15460
rect 13202 15307 13212 15460
rect 13278 15307 13288 15460
rect 13394 15307 13404 15460
rect 13470 15307 13480 15460
rect 13586 15307 13596 15460
rect 13662 15307 13672 15460
rect 13778 15307 13788 15460
rect 13854 15307 13864 15460
rect 13970 15307 13980 15460
rect 14046 15307 14056 15460
rect 14162 15307 14172 15460
rect 14238 15307 14248 15460
rect 14284 15247 14504 15494
rect 14646 15307 14656 15460
rect 14722 15307 14732 15460
rect 14838 15307 14848 15460
rect 14914 15307 14924 15460
rect 15030 15307 15040 15460
rect 15106 15307 15116 15460
rect 15222 15307 15232 15460
rect 15298 15307 15308 15460
rect 15414 15307 15424 15460
rect 15490 15307 15500 15460
rect 15606 15307 15616 15460
rect 15682 15307 15692 15460
rect 15798 15307 15808 15460
rect 15874 15307 15884 15460
rect 15990 15307 16000 15460
rect 16066 15307 16076 15460
rect 16112 15247 16332 15494
rect 16474 15307 16484 15460
rect 16550 15307 16560 15460
rect 16666 15307 16676 15460
rect 16742 15307 16752 15460
rect 16858 15307 16868 15460
rect 16934 15307 16944 15460
rect 17050 15307 17060 15460
rect 17126 15307 17136 15460
rect 17242 15307 17252 15460
rect 17318 15307 17328 15460
rect 17434 15307 17444 15460
rect 17510 15307 17520 15460
rect 17626 15307 17636 15460
rect 17702 15307 17712 15460
rect 17818 15307 17828 15460
rect 17894 15307 17904 15460
rect 17940 15247 18160 15494
rect 18302 15307 18312 15460
rect 18378 15307 18388 15460
rect 18494 15307 18504 15460
rect 18570 15307 18580 15460
rect 18686 15307 18696 15460
rect 18762 15307 18772 15460
rect 18878 15307 18888 15460
rect 18954 15307 18964 15460
rect 19070 15307 19080 15460
rect 19146 15307 19156 15460
rect 19262 15307 19272 15460
rect 19338 15307 19348 15460
rect 19454 15307 19464 15460
rect 19530 15307 19540 15460
rect 19646 15307 19656 15460
rect 19722 15307 19732 15460
rect 19768 15247 19988 15494
rect 20130 15307 20140 15460
rect 20206 15307 20216 15460
rect 20322 15307 20332 15460
rect 20398 15307 20408 15460
rect 20514 15307 20524 15460
rect 20590 15307 20600 15460
rect 20706 15307 20716 15460
rect 20782 15307 20792 15460
rect 20898 15307 20908 15460
rect 20974 15307 20984 15460
rect 21090 15307 21100 15460
rect 21166 15307 21176 15460
rect 21282 15307 21292 15460
rect 21358 15307 21368 15460
rect 21474 15307 21484 15460
rect 21550 15307 21560 15460
rect 21596 15247 21816 15494
rect 118 15094 128 15247
rect 194 15094 204 15247
rect 310 15094 320 15247
rect 386 15094 396 15247
rect 502 15094 512 15247
rect 578 15094 588 15247
rect 694 15094 704 15247
rect 770 15094 780 15247
rect 886 15094 896 15247
rect 962 15094 972 15247
rect 1078 15094 1088 15247
rect 1154 15094 1164 15247
rect 1270 15094 1280 15247
rect 1346 15094 1356 15247
rect 1462 15094 1472 15247
rect 1528 15094 1708 15247
rect 1946 15094 1956 15247
rect 2022 15094 2032 15247
rect 2138 15094 2148 15247
rect 2214 15094 2224 15247
rect 2330 15094 2340 15247
rect 2406 15094 2416 15247
rect 2522 15094 2532 15247
rect 2598 15094 2608 15247
rect 2714 15094 2724 15247
rect 2790 15094 2800 15247
rect 2906 15094 2916 15247
rect 2982 15094 2992 15247
rect 3098 15094 3108 15247
rect 3174 15094 3184 15247
rect 3290 15094 3300 15247
rect 3356 15094 3536 15247
rect 3774 15094 3784 15247
rect 3850 15094 3860 15247
rect 3966 15094 3976 15247
rect 4042 15094 4052 15247
rect 4158 15094 4168 15247
rect 4234 15094 4244 15247
rect 4350 15094 4360 15247
rect 4426 15094 4436 15247
rect 4542 15094 4552 15247
rect 4618 15094 4628 15247
rect 4734 15094 4744 15247
rect 4810 15094 4820 15247
rect 4926 15094 4936 15247
rect 5002 15094 5012 15247
rect 5118 15094 5128 15247
rect 5184 15094 5364 15247
rect 5602 15094 5612 15247
rect 5678 15094 5688 15247
rect 5794 15094 5804 15247
rect 5870 15094 5880 15247
rect 5986 15094 5996 15247
rect 6062 15094 6072 15247
rect 6178 15094 6188 15247
rect 6254 15094 6264 15247
rect 6370 15094 6380 15247
rect 6446 15094 6456 15247
rect 6562 15094 6572 15247
rect 6638 15094 6648 15247
rect 6754 15094 6764 15247
rect 6830 15094 6840 15247
rect 6946 15094 6956 15247
rect 7012 15094 7192 15247
rect 7430 15094 7440 15247
rect 7506 15094 7516 15247
rect 7622 15094 7632 15247
rect 7698 15094 7708 15247
rect 7814 15094 7824 15247
rect 7890 15094 7900 15247
rect 8006 15094 8016 15247
rect 8082 15094 8092 15247
rect 8198 15094 8208 15247
rect 8274 15094 8284 15247
rect 8390 15094 8400 15247
rect 8466 15094 8476 15247
rect 8582 15094 8592 15247
rect 8658 15094 8668 15247
rect 8774 15094 8784 15247
rect 8840 15094 9020 15247
rect 9258 15094 9268 15247
rect 9334 15094 9344 15247
rect 9450 15094 9460 15247
rect 9526 15094 9536 15247
rect 9642 15094 9652 15247
rect 9718 15094 9728 15247
rect 9834 15094 9844 15247
rect 9910 15094 9920 15247
rect 10026 15094 10036 15247
rect 10102 15094 10112 15247
rect 10218 15094 10228 15247
rect 10294 15094 10304 15247
rect 10410 15094 10420 15247
rect 10486 15094 10496 15247
rect 10602 15094 10612 15247
rect 10668 15094 10848 15247
rect 11086 15094 11096 15247
rect 11162 15094 11172 15247
rect 11278 15094 11288 15247
rect 11354 15094 11364 15247
rect 11470 15094 11480 15247
rect 11546 15094 11556 15247
rect 11662 15094 11672 15247
rect 11738 15094 11748 15247
rect 11854 15094 11864 15247
rect 11930 15094 11940 15247
rect 12046 15094 12056 15247
rect 12122 15094 12132 15247
rect 12238 15094 12248 15247
rect 12314 15094 12324 15247
rect 12430 15094 12440 15247
rect 12496 15094 12676 15247
rect 12914 15094 12924 15247
rect 12990 15094 13000 15247
rect 13106 15094 13116 15247
rect 13182 15094 13192 15247
rect 13298 15094 13308 15247
rect 13374 15094 13384 15247
rect 13490 15094 13500 15247
rect 13566 15094 13576 15247
rect 13682 15094 13692 15247
rect 13758 15094 13768 15247
rect 13874 15094 13884 15247
rect 13950 15094 13960 15247
rect 14066 15094 14076 15247
rect 14142 15094 14152 15247
rect 14258 15094 14268 15247
rect 14324 15094 14504 15247
rect 14742 15094 14752 15247
rect 14818 15094 14828 15247
rect 14934 15094 14944 15247
rect 15010 15094 15020 15247
rect 15126 15094 15136 15247
rect 15202 15094 15212 15247
rect 15318 15094 15328 15247
rect 15394 15094 15404 15247
rect 15510 15094 15520 15247
rect 15586 15094 15596 15247
rect 15702 15094 15712 15247
rect 15778 15094 15788 15247
rect 15894 15094 15904 15247
rect 15970 15094 15980 15247
rect 16086 15094 16096 15247
rect 16152 15094 16332 15247
rect 16570 15094 16580 15247
rect 16646 15094 16656 15247
rect 16762 15094 16772 15247
rect 16838 15094 16848 15247
rect 16954 15094 16964 15247
rect 17030 15094 17040 15247
rect 17146 15094 17156 15247
rect 17222 15094 17232 15247
rect 17338 15094 17348 15247
rect 17414 15094 17424 15247
rect 17530 15094 17540 15247
rect 17606 15094 17616 15247
rect 17722 15094 17732 15247
rect 17798 15094 17808 15247
rect 17914 15094 17924 15247
rect 17980 15094 18160 15247
rect 18398 15094 18408 15247
rect 18474 15094 18484 15247
rect 18590 15094 18600 15247
rect 18666 15094 18676 15247
rect 18782 15094 18792 15247
rect 18858 15094 18868 15247
rect 18974 15094 18984 15247
rect 19050 15094 19060 15247
rect 19166 15094 19176 15247
rect 19242 15094 19252 15247
rect 19358 15094 19368 15247
rect 19434 15094 19444 15247
rect 19550 15094 19560 15247
rect 19626 15094 19636 15247
rect 19742 15094 19752 15247
rect 19808 15094 19988 15247
rect 20226 15094 20236 15247
rect 20302 15094 20312 15247
rect 20418 15094 20428 15247
rect 20494 15094 20504 15247
rect 20610 15094 20620 15247
rect 20686 15094 20696 15247
rect 20802 15094 20812 15247
rect 20878 15094 20888 15247
rect 20994 15094 21004 15247
rect 21070 15094 21080 15247
rect 21186 15094 21196 15247
rect 21262 15094 21272 15247
rect 21378 15094 21388 15247
rect 21454 15094 21464 15247
rect 21570 15094 21580 15247
rect 21636 15094 21816 15247
rect 0 14997 1490 15056
rect 1828 14997 3318 15056
rect 3656 14997 5146 15056
rect 5484 14997 6974 15056
rect 7312 14997 8802 15056
rect 9140 14997 10630 15056
rect 10968 14997 12458 15056
rect 12796 14997 14286 15056
rect 14624 14997 16114 15056
rect 16452 14997 17942 15056
rect 18280 14997 19770 15056
rect 20108 14997 21598 15056
rect 0 14818 1490 14877
rect 1828 14818 3318 14877
rect 3656 14818 5146 14877
rect 5484 14818 6974 14877
rect 7312 14818 8802 14877
rect 9140 14818 10630 14877
rect 10968 14818 12458 14877
rect 12796 14818 14286 14877
rect 14624 14818 16114 14877
rect 16452 14818 17942 14877
rect 18280 14818 19770 14877
rect 20108 14818 21598 14877
rect 22 14593 32 14746
rect 98 14593 108 14746
rect 214 14593 224 14746
rect 290 14593 300 14746
rect 406 14593 416 14746
rect 482 14593 492 14746
rect 598 14593 608 14746
rect 674 14593 684 14746
rect 790 14593 800 14746
rect 866 14593 876 14746
rect 982 14593 992 14746
rect 1058 14593 1068 14746
rect 1174 14593 1184 14746
rect 1250 14593 1260 14746
rect 1366 14593 1376 14746
rect 1442 14593 1452 14746
rect 1488 14533 1708 14780
rect 1850 14593 1860 14746
rect 1926 14593 1936 14746
rect 2042 14593 2052 14746
rect 2118 14593 2128 14746
rect 2234 14593 2244 14746
rect 2310 14593 2320 14746
rect 2426 14593 2436 14746
rect 2502 14593 2512 14746
rect 2618 14593 2628 14746
rect 2694 14593 2704 14746
rect 2810 14593 2820 14746
rect 2886 14593 2896 14746
rect 3002 14593 3012 14746
rect 3078 14593 3088 14746
rect 3194 14593 3204 14746
rect 3270 14593 3280 14746
rect 3316 14533 3536 14780
rect 3678 14593 3688 14746
rect 3754 14593 3764 14746
rect 3870 14593 3880 14746
rect 3946 14593 3956 14746
rect 4062 14593 4072 14746
rect 4138 14593 4148 14746
rect 4254 14593 4264 14746
rect 4330 14593 4340 14746
rect 4446 14593 4456 14746
rect 4522 14593 4532 14746
rect 4638 14593 4648 14746
rect 4714 14593 4724 14746
rect 4830 14593 4840 14746
rect 4906 14593 4916 14746
rect 5022 14593 5032 14746
rect 5098 14593 5108 14746
rect 5144 14533 5364 14780
rect 5506 14593 5516 14746
rect 5582 14593 5592 14746
rect 5698 14593 5708 14746
rect 5774 14593 5784 14746
rect 5890 14593 5900 14746
rect 5966 14593 5976 14746
rect 6082 14593 6092 14746
rect 6158 14593 6168 14746
rect 6274 14593 6284 14746
rect 6350 14593 6360 14746
rect 6466 14593 6476 14746
rect 6542 14593 6552 14746
rect 6658 14593 6668 14746
rect 6734 14593 6744 14746
rect 6850 14593 6860 14746
rect 6926 14593 6936 14746
rect 6972 14533 7192 14780
rect 7334 14593 7344 14746
rect 7410 14593 7420 14746
rect 7526 14593 7536 14746
rect 7602 14593 7612 14746
rect 7718 14593 7728 14746
rect 7794 14593 7804 14746
rect 7910 14593 7920 14746
rect 7986 14593 7996 14746
rect 8102 14593 8112 14746
rect 8178 14593 8188 14746
rect 8294 14593 8304 14746
rect 8370 14593 8380 14746
rect 8486 14593 8496 14746
rect 8562 14593 8572 14746
rect 8678 14593 8688 14746
rect 8754 14593 8764 14746
rect 8800 14533 9020 14780
rect 9162 14593 9172 14746
rect 9238 14593 9248 14746
rect 9354 14593 9364 14746
rect 9430 14593 9440 14746
rect 9546 14593 9556 14746
rect 9622 14593 9632 14746
rect 9738 14593 9748 14746
rect 9814 14593 9824 14746
rect 9930 14593 9940 14746
rect 10006 14593 10016 14746
rect 10122 14593 10132 14746
rect 10198 14593 10208 14746
rect 10314 14593 10324 14746
rect 10390 14593 10400 14746
rect 10506 14593 10516 14746
rect 10582 14593 10592 14746
rect 10628 14533 10848 14780
rect 10990 14593 11000 14746
rect 11066 14593 11076 14746
rect 11182 14593 11192 14746
rect 11258 14593 11268 14746
rect 11374 14593 11384 14746
rect 11450 14593 11460 14746
rect 11566 14593 11576 14746
rect 11642 14593 11652 14746
rect 11758 14593 11768 14746
rect 11834 14593 11844 14746
rect 11950 14593 11960 14746
rect 12026 14593 12036 14746
rect 12142 14593 12152 14746
rect 12218 14593 12228 14746
rect 12334 14593 12344 14746
rect 12410 14593 12420 14746
rect 12456 14533 12676 14780
rect 12818 14593 12828 14746
rect 12894 14593 12904 14746
rect 13010 14593 13020 14746
rect 13086 14593 13096 14746
rect 13202 14593 13212 14746
rect 13278 14593 13288 14746
rect 13394 14593 13404 14746
rect 13470 14593 13480 14746
rect 13586 14593 13596 14746
rect 13662 14593 13672 14746
rect 13778 14593 13788 14746
rect 13854 14593 13864 14746
rect 13970 14593 13980 14746
rect 14046 14593 14056 14746
rect 14162 14593 14172 14746
rect 14238 14593 14248 14746
rect 14284 14533 14504 14780
rect 14646 14593 14656 14746
rect 14722 14593 14732 14746
rect 14838 14593 14848 14746
rect 14914 14593 14924 14746
rect 15030 14593 15040 14746
rect 15106 14593 15116 14746
rect 15222 14593 15232 14746
rect 15298 14593 15308 14746
rect 15414 14593 15424 14746
rect 15490 14593 15500 14746
rect 15606 14593 15616 14746
rect 15682 14593 15692 14746
rect 15798 14593 15808 14746
rect 15874 14593 15884 14746
rect 15990 14593 16000 14746
rect 16066 14593 16076 14746
rect 16112 14533 16332 14780
rect 16474 14593 16484 14746
rect 16550 14593 16560 14746
rect 16666 14593 16676 14746
rect 16742 14593 16752 14746
rect 16858 14593 16868 14746
rect 16934 14593 16944 14746
rect 17050 14593 17060 14746
rect 17126 14593 17136 14746
rect 17242 14593 17252 14746
rect 17318 14593 17328 14746
rect 17434 14593 17444 14746
rect 17510 14593 17520 14746
rect 17626 14593 17636 14746
rect 17702 14593 17712 14746
rect 17818 14593 17828 14746
rect 17894 14593 17904 14746
rect 17940 14533 18160 14780
rect 18302 14593 18312 14746
rect 18378 14593 18388 14746
rect 18494 14593 18504 14746
rect 18570 14593 18580 14746
rect 18686 14593 18696 14746
rect 18762 14593 18772 14746
rect 18878 14593 18888 14746
rect 18954 14593 18964 14746
rect 19070 14593 19080 14746
rect 19146 14593 19156 14746
rect 19262 14593 19272 14746
rect 19338 14593 19348 14746
rect 19454 14593 19464 14746
rect 19530 14593 19540 14746
rect 19646 14593 19656 14746
rect 19722 14593 19732 14746
rect 19768 14533 19988 14780
rect 20130 14593 20140 14746
rect 20206 14593 20216 14746
rect 20322 14593 20332 14746
rect 20398 14593 20408 14746
rect 20514 14593 20524 14746
rect 20590 14593 20600 14746
rect 20706 14593 20716 14746
rect 20782 14593 20792 14746
rect 20898 14593 20908 14746
rect 20974 14593 20984 14746
rect 21090 14593 21100 14746
rect 21166 14593 21176 14746
rect 21282 14593 21292 14746
rect 21358 14593 21368 14746
rect 21474 14593 21484 14746
rect 21550 14593 21560 14746
rect 21596 14533 21816 14780
rect 118 14380 128 14533
rect 194 14380 204 14533
rect 310 14380 320 14533
rect 386 14380 396 14533
rect 502 14380 512 14533
rect 578 14380 588 14533
rect 694 14380 704 14533
rect 770 14380 780 14533
rect 886 14380 896 14533
rect 962 14380 972 14533
rect 1078 14380 1088 14533
rect 1154 14380 1164 14533
rect 1270 14380 1280 14533
rect 1346 14380 1356 14533
rect 1462 14380 1472 14533
rect 1528 14380 1708 14533
rect 1946 14380 1956 14533
rect 2022 14380 2032 14533
rect 2138 14380 2148 14533
rect 2214 14380 2224 14533
rect 2330 14380 2340 14533
rect 2406 14380 2416 14533
rect 2522 14380 2532 14533
rect 2598 14380 2608 14533
rect 2714 14380 2724 14533
rect 2790 14380 2800 14533
rect 2906 14380 2916 14533
rect 2982 14380 2992 14533
rect 3098 14380 3108 14533
rect 3174 14380 3184 14533
rect 3290 14380 3300 14533
rect 3356 14380 3536 14533
rect 3774 14380 3784 14533
rect 3850 14380 3860 14533
rect 3966 14380 3976 14533
rect 4042 14380 4052 14533
rect 4158 14380 4168 14533
rect 4234 14380 4244 14533
rect 4350 14380 4360 14533
rect 4426 14380 4436 14533
rect 4542 14380 4552 14533
rect 4618 14380 4628 14533
rect 4734 14380 4744 14533
rect 4810 14380 4820 14533
rect 4926 14380 4936 14533
rect 5002 14380 5012 14533
rect 5118 14380 5128 14533
rect 5184 14380 5364 14533
rect 5602 14380 5612 14533
rect 5678 14380 5688 14533
rect 5794 14380 5804 14533
rect 5870 14380 5880 14533
rect 5986 14380 5996 14533
rect 6062 14380 6072 14533
rect 6178 14380 6188 14533
rect 6254 14380 6264 14533
rect 6370 14380 6380 14533
rect 6446 14380 6456 14533
rect 6562 14380 6572 14533
rect 6638 14380 6648 14533
rect 6754 14380 6764 14533
rect 6830 14380 6840 14533
rect 6946 14380 6956 14533
rect 7012 14380 7192 14533
rect 7430 14380 7440 14533
rect 7506 14380 7516 14533
rect 7622 14380 7632 14533
rect 7698 14380 7708 14533
rect 7814 14380 7824 14533
rect 7890 14380 7900 14533
rect 8006 14380 8016 14533
rect 8082 14380 8092 14533
rect 8198 14380 8208 14533
rect 8274 14380 8284 14533
rect 8390 14380 8400 14533
rect 8466 14380 8476 14533
rect 8582 14380 8592 14533
rect 8658 14380 8668 14533
rect 8774 14380 8784 14533
rect 8840 14380 9020 14533
rect 9258 14380 9268 14533
rect 9334 14380 9344 14533
rect 9450 14380 9460 14533
rect 9526 14380 9536 14533
rect 9642 14380 9652 14533
rect 9718 14380 9728 14533
rect 9834 14380 9844 14533
rect 9910 14380 9920 14533
rect 10026 14380 10036 14533
rect 10102 14380 10112 14533
rect 10218 14380 10228 14533
rect 10294 14380 10304 14533
rect 10410 14380 10420 14533
rect 10486 14380 10496 14533
rect 10602 14380 10612 14533
rect 10668 14380 10848 14533
rect 11086 14380 11096 14533
rect 11162 14380 11172 14533
rect 11278 14380 11288 14533
rect 11354 14380 11364 14533
rect 11470 14380 11480 14533
rect 11546 14380 11556 14533
rect 11662 14380 11672 14533
rect 11738 14380 11748 14533
rect 11854 14380 11864 14533
rect 11930 14380 11940 14533
rect 12046 14380 12056 14533
rect 12122 14380 12132 14533
rect 12238 14380 12248 14533
rect 12314 14380 12324 14533
rect 12430 14380 12440 14533
rect 12496 14380 12676 14533
rect 12914 14380 12924 14533
rect 12990 14380 13000 14533
rect 13106 14380 13116 14533
rect 13182 14380 13192 14533
rect 13298 14380 13308 14533
rect 13374 14380 13384 14533
rect 13490 14380 13500 14533
rect 13566 14380 13576 14533
rect 13682 14380 13692 14533
rect 13758 14380 13768 14533
rect 13874 14380 13884 14533
rect 13950 14380 13960 14533
rect 14066 14380 14076 14533
rect 14142 14380 14152 14533
rect 14258 14380 14268 14533
rect 14324 14380 14504 14533
rect 14742 14380 14752 14533
rect 14818 14380 14828 14533
rect 14934 14380 14944 14533
rect 15010 14380 15020 14533
rect 15126 14380 15136 14533
rect 15202 14380 15212 14533
rect 15318 14380 15328 14533
rect 15394 14380 15404 14533
rect 15510 14380 15520 14533
rect 15586 14380 15596 14533
rect 15702 14380 15712 14533
rect 15778 14380 15788 14533
rect 15894 14380 15904 14533
rect 15970 14380 15980 14533
rect 16086 14380 16096 14533
rect 16152 14380 16332 14533
rect 16570 14380 16580 14533
rect 16646 14380 16656 14533
rect 16762 14380 16772 14533
rect 16838 14380 16848 14533
rect 16954 14380 16964 14533
rect 17030 14380 17040 14533
rect 17146 14380 17156 14533
rect 17222 14380 17232 14533
rect 17338 14380 17348 14533
rect 17414 14380 17424 14533
rect 17530 14380 17540 14533
rect 17606 14380 17616 14533
rect 17722 14380 17732 14533
rect 17798 14380 17808 14533
rect 17914 14380 17924 14533
rect 17980 14380 18160 14533
rect 18398 14380 18408 14533
rect 18474 14380 18484 14533
rect 18590 14380 18600 14533
rect 18666 14380 18676 14533
rect 18782 14380 18792 14533
rect 18858 14380 18868 14533
rect 18974 14380 18984 14533
rect 19050 14380 19060 14533
rect 19166 14380 19176 14533
rect 19242 14380 19252 14533
rect 19358 14380 19368 14533
rect 19434 14380 19444 14533
rect 19550 14380 19560 14533
rect 19626 14380 19636 14533
rect 19742 14380 19752 14533
rect 19808 14380 19988 14533
rect 20226 14380 20236 14533
rect 20302 14380 20312 14533
rect 20418 14380 20428 14533
rect 20494 14380 20504 14533
rect 20610 14380 20620 14533
rect 20686 14380 20696 14533
rect 20802 14380 20812 14533
rect 20878 14380 20888 14533
rect 20994 14380 21004 14533
rect 21070 14380 21080 14533
rect 21186 14380 21196 14533
rect 21262 14380 21272 14533
rect 21378 14380 21388 14533
rect 21454 14380 21464 14533
rect 21570 14380 21580 14533
rect 21636 14380 21816 14533
rect 0 14283 1490 14342
rect 1828 14283 3318 14342
rect 3656 14283 5146 14342
rect 5484 14283 6974 14342
rect 7312 14283 8802 14342
rect 9140 14283 10630 14342
rect 10968 14283 12458 14342
rect 12796 14283 14286 14342
rect 14624 14283 16114 14342
rect 16452 14283 17942 14342
rect 18280 14283 19770 14342
rect 20108 14283 21598 14342
rect 0 14104 1490 14163
rect 1828 14104 3318 14163
rect 3656 14104 5146 14163
rect 5484 14104 6974 14163
rect 7312 14104 8802 14163
rect 9140 14104 10630 14163
rect 10968 14104 12458 14163
rect 12796 14104 14286 14163
rect 14624 14104 16114 14163
rect 16452 14104 17942 14163
rect 18280 14104 19770 14163
rect 20108 14104 21598 14163
rect 22 13879 32 14032
rect 98 13879 108 14032
rect 214 13879 224 14032
rect 290 13879 300 14032
rect 406 13879 416 14032
rect 482 13879 492 14032
rect 598 13879 608 14032
rect 674 13879 684 14032
rect 790 13879 800 14032
rect 866 13879 876 14032
rect 982 13879 992 14032
rect 1058 13879 1068 14032
rect 1174 13879 1184 14032
rect 1250 13879 1260 14032
rect 1366 13879 1376 14032
rect 1442 13879 1452 14032
rect 1488 13819 1708 14066
rect 1850 13879 1860 14032
rect 1926 13879 1936 14032
rect 2042 13879 2052 14032
rect 2118 13879 2128 14032
rect 2234 13879 2244 14032
rect 2310 13879 2320 14032
rect 2426 13879 2436 14032
rect 2502 13879 2512 14032
rect 2618 13879 2628 14032
rect 2694 13879 2704 14032
rect 2810 13879 2820 14032
rect 2886 13879 2896 14032
rect 3002 13879 3012 14032
rect 3078 13879 3088 14032
rect 3194 13879 3204 14032
rect 3270 13879 3280 14032
rect 3316 13819 3536 14066
rect 3678 13879 3688 14032
rect 3754 13879 3764 14032
rect 3870 13879 3880 14032
rect 3946 13879 3956 14032
rect 4062 13879 4072 14032
rect 4138 13879 4148 14032
rect 4254 13879 4264 14032
rect 4330 13879 4340 14032
rect 4446 13879 4456 14032
rect 4522 13879 4532 14032
rect 4638 13879 4648 14032
rect 4714 13879 4724 14032
rect 4830 13879 4840 14032
rect 4906 13879 4916 14032
rect 5022 13879 5032 14032
rect 5098 13879 5108 14032
rect 5144 13819 5364 14066
rect 5506 13879 5516 14032
rect 5582 13879 5592 14032
rect 5698 13879 5708 14032
rect 5774 13879 5784 14032
rect 5890 13879 5900 14032
rect 5966 13879 5976 14032
rect 6082 13879 6092 14032
rect 6158 13879 6168 14032
rect 6274 13879 6284 14032
rect 6350 13879 6360 14032
rect 6466 13879 6476 14032
rect 6542 13879 6552 14032
rect 6658 13879 6668 14032
rect 6734 13879 6744 14032
rect 6850 13879 6860 14032
rect 6926 13879 6936 14032
rect 6972 13819 7192 14066
rect 7334 13879 7344 14032
rect 7410 13879 7420 14032
rect 7526 13879 7536 14032
rect 7602 13879 7612 14032
rect 7718 13879 7728 14032
rect 7794 13879 7804 14032
rect 7910 13879 7920 14032
rect 7986 13879 7996 14032
rect 8102 13879 8112 14032
rect 8178 13879 8188 14032
rect 8294 13879 8304 14032
rect 8370 13879 8380 14032
rect 8486 13879 8496 14032
rect 8562 13879 8572 14032
rect 8678 13879 8688 14032
rect 8754 13879 8764 14032
rect 8800 13819 9020 14066
rect 9162 13879 9172 14032
rect 9238 13879 9248 14032
rect 9354 13879 9364 14032
rect 9430 13879 9440 14032
rect 9546 13879 9556 14032
rect 9622 13879 9632 14032
rect 9738 13879 9748 14032
rect 9814 13879 9824 14032
rect 9930 13879 9940 14032
rect 10006 13879 10016 14032
rect 10122 13879 10132 14032
rect 10198 13879 10208 14032
rect 10314 13879 10324 14032
rect 10390 13879 10400 14032
rect 10506 13879 10516 14032
rect 10582 13879 10592 14032
rect 10628 13819 10848 14066
rect 10990 13879 11000 14032
rect 11066 13879 11076 14032
rect 11182 13879 11192 14032
rect 11258 13879 11268 14032
rect 11374 13879 11384 14032
rect 11450 13879 11460 14032
rect 11566 13879 11576 14032
rect 11642 13879 11652 14032
rect 11758 13879 11768 14032
rect 11834 13879 11844 14032
rect 11950 13879 11960 14032
rect 12026 13879 12036 14032
rect 12142 13879 12152 14032
rect 12218 13879 12228 14032
rect 12334 13879 12344 14032
rect 12410 13879 12420 14032
rect 12456 13819 12676 14066
rect 12818 13879 12828 14032
rect 12894 13879 12904 14032
rect 13010 13879 13020 14032
rect 13086 13879 13096 14032
rect 13202 13879 13212 14032
rect 13278 13879 13288 14032
rect 13394 13879 13404 14032
rect 13470 13879 13480 14032
rect 13586 13879 13596 14032
rect 13662 13879 13672 14032
rect 13778 13879 13788 14032
rect 13854 13879 13864 14032
rect 13970 13879 13980 14032
rect 14046 13879 14056 14032
rect 14162 13879 14172 14032
rect 14238 13879 14248 14032
rect 14284 13819 14504 14066
rect 14646 13879 14656 14032
rect 14722 13879 14732 14032
rect 14838 13879 14848 14032
rect 14914 13879 14924 14032
rect 15030 13879 15040 14032
rect 15106 13879 15116 14032
rect 15222 13879 15232 14032
rect 15298 13879 15308 14032
rect 15414 13879 15424 14032
rect 15490 13879 15500 14032
rect 15606 13879 15616 14032
rect 15682 13879 15692 14032
rect 15798 13879 15808 14032
rect 15874 13879 15884 14032
rect 15990 13879 16000 14032
rect 16066 13879 16076 14032
rect 16112 13819 16332 14066
rect 16474 13879 16484 14032
rect 16550 13879 16560 14032
rect 16666 13879 16676 14032
rect 16742 13879 16752 14032
rect 16858 13879 16868 14032
rect 16934 13879 16944 14032
rect 17050 13879 17060 14032
rect 17126 13879 17136 14032
rect 17242 13879 17252 14032
rect 17318 13879 17328 14032
rect 17434 13879 17444 14032
rect 17510 13879 17520 14032
rect 17626 13879 17636 14032
rect 17702 13879 17712 14032
rect 17818 13879 17828 14032
rect 17894 13879 17904 14032
rect 17940 13819 18160 14066
rect 18302 13879 18312 14032
rect 18378 13879 18388 14032
rect 18494 13879 18504 14032
rect 18570 13879 18580 14032
rect 18686 13879 18696 14032
rect 18762 13879 18772 14032
rect 18878 13879 18888 14032
rect 18954 13879 18964 14032
rect 19070 13879 19080 14032
rect 19146 13879 19156 14032
rect 19262 13879 19272 14032
rect 19338 13879 19348 14032
rect 19454 13879 19464 14032
rect 19530 13879 19540 14032
rect 19646 13879 19656 14032
rect 19722 13879 19732 14032
rect 19768 13819 19988 14066
rect 20130 13879 20140 14032
rect 20206 13879 20216 14032
rect 20322 13879 20332 14032
rect 20398 13879 20408 14032
rect 20514 13879 20524 14032
rect 20590 13879 20600 14032
rect 20706 13879 20716 14032
rect 20782 13879 20792 14032
rect 20898 13879 20908 14032
rect 20974 13879 20984 14032
rect 21090 13879 21100 14032
rect 21166 13879 21176 14032
rect 21282 13879 21292 14032
rect 21358 13879 21368 14032
rect 21474 13879 21484 14032
rect 21550 13879 21560 14032
rect 21596 13819 21816 14066
rect 118 13666 128 13819
rect 194 13666 204 13819
rect 310 13666 320 13819
rect 386 13666 396 13819
rect 502 13666 512 13819
rect 578 13666 588 13819
rect 694 13666 704 13819
rect 770 13666 780 13819
rect 886 13666 896 13819
rect 962 13666 972 13819
rect 1078 13666 1088 13819
rect 1154 13666 1164 13819
rect 1270 13666 1280 13819
rect 1346 13666 1356 13819
rect 1462 13666 1472 13819
rect 1528 13666 1708 13819
rect 1946 13666 1956 13819
rect 2022 13666 2032 13819
rect 2138 13666 2148 13819
rect 2214 13666 2224 13819
rect 2330 13666 2340 13819
rect 2406 13666 2416 13819
rect 2522 13666 2532 13819
rect 2598 13666 2608 13819
rect 2714 13666 2724 13819
rect 2790 13666 2800 13819
rect 2906 13666 2916 13819
rect 2982 13666 2992 13819
rect 3098 13666 3108 13819
rect 3174 13666 3184 13819
rect 3290 13666 3300 13819
rect 3356 13666 3536 13819
rect 3774 13666 3784 13819
rect 3850 13666 3860 13819
rect 3966 13666 3976 13819
rect 4042 13666 4052 13819
rect 4158 13666 4168 13819
rect 4234 13666 4244 13819
rect 4350 13666 4360 13819
rect 4426 13666 4436 13819
rect 4542 13666 4552 13819
rect 4618 13666 4628 13819
rect 4734 13666 4744 13819
rect 4810 13666 4820 13819
rect 4926 13666 4936 13819
rect 5002 13666 5012 13819
rect 5118 13666 5128 13819
rect 5184 13666 5364 13819
rect 5602 13666 5612 13819
rect 5678 13666 5688 13819
rect 5794 13666 5804 13819
rect 5870 13666 5880 13819
rect 5986 13666 5996 13819
rect 6062 13666 6072 13819
rect 6178 13666 6188 13819
rect 6254 13666 6264 13819
rect 6370 13666 6380 13819
rect 6446 13666 6456 13819
rect 6562 13666 6572 13819
rect 6638 13666 6648 13819
rect 6754 13666 6764 13819
rect 6830 13666 6840 13819
rect 6946 13666 6956 13819
rect 7012 13666 7192 13819
rect 7430 13666 7440 13819
rect 7506 13666 7516 13819
rect 7622 13666 7632 13819
rect 7698 13666 7708 13819
rect 7814 13666 7824 13819
rect 7890 13666 7900 13819
rect 8006 13666 8016 13819
rect 8082 13666 8092 13819
rect 8198 13666 8208 13819
rect 8274 13666 8284 13819
rect 8390 13666 8400 13819
rect 8466 13666 8476 13819
rect 8582 13666 8592 13819
rect 8658 13666 8668 13819
rect 8774 13666 8784 13819
rect 8840 13666 9020 13819
rect 9258 13666 9268 13819
rect 9334 13666 9344 13819
rect 9450 13666 9460 13819
rect 9526 13666 9536 13819
rect 9642 13666 9652 13819
rect 9718 13666 9728 13819
rect 9834 13666 9844 13819
rect 9910 13666 9920 13819
rect 10026 13666 10036 13819
rect 10102 13666 10112 13819
rect 10218 13666 10228 13819
rect 10294 13666 10304 13819
rect 10410 13666 10420 13819
rect 10486 13666 10496 13819
rect 10602 13666 10612 13819
rect 10668 13666 10848 13819
rect 11086 13666 11096 13819
rect 11162 13666 11172 13819
rect 11278 13666 11288 13819
rect 11354 13666 11364 13819
rect 11470 13666 11480 13819
rect 11546 13666 11556 13819
rect 11662 13666 11672 13819
rect 11738 13666 11748 13819
rect 11854 13666 11864 13819
rect 11930 13666 11940 13819
rect 12046 13666 12056 13819
rect 12122 13666 12132 13819
rect 12238 13666 12248 13819
rect 12314 13666 12324 13819
rect 12430 13666 12440 13819
rect 12496 13666 12676 13819
rect 12914 13666 12924 13819
rect 12990 13666 13000 13819
rect 13106 13666 13116 13819
rect 13182 13666 13192 13819
rect 13298 13666 13308 13819
rect 13374 13666 13384 13819
rect 13490 13666 13500 13819
rect 13566 13666 13576 13819
rect 13682 13666 13692 13819
rect 13758 13666 13768 13819
rect 13874 13666 13884 13819
rect 13950 13666 13960 13819
rect 14066 13666 14076 13819
rect 14142 13666 14152 13819
rect 14258 13666 14268 13819
rect 14324 13666 14504 13819
rect 14742 13666 14752 13819
rect 14818 13666 14828 13819
rect 14934 13666 14944 13819
rect 15010 13666 15020 13819
rect 15126 13666 15136 13819
rect 15202 13666 15212 13819
rect 15318 13666 15328 13819
rect 15394 13666 15404 13819
rect 15510 13666 15520 13819
rect 15586 13666 15596 13819
rect 15702 13666 15712 13819
rect 15778 13666 15788 13819
rect 15894 13666 15904 13819
rect 15970 13666 15980 13819
rect 16086 13666 16096 13819
rect 16152 13666 16332 13819
rect 16570 13666 16580 13819
rect 16646 13666 16656 13819
rect 16762 13666 16772 13819
rect 16838 13666 16848 13819
rect 16954 13666 16964 13819
rect 17030 13666 17040 13819
rect 17146 13666 17156 13819
rect 17222 13666 17232 13819
rect 17338 13666 17348 13819
rect 17414 13666 17424 13819
rect 17530 13666 17540 13819
rect 17606 13666 17616 13819
rect 17722 13666 17732 13819
rect 17798 13666 17808 13819
rect 17914 13666 17924 13819
rect 17980 13666 18160 13819
rect 18398 13666 18408 13819
rect 18474 13666 18484 13819
rect 18590 13666 18600 13819
rect 18666 13666 18676 13819
rect 18782 13666 18792 13819
rect 18858 13666 18868 13819
rect 18974 13666 18984 13819
rect 19050 13666 19060 13819
rect 19166 13666 19176 13819
rect 19242 13666 19252 13819
rect 19358 13666 19368 13819
rect 19434 13666 19444 13819
rect 19550 13666 19560 13819
rect 19626 13666 19636 13819
rect 19742 13666 19752 13819
rect 19808 13666 19988 13819
rect 20226 13666 20236 13819
rect 20302 13666 20312 13819
rect 20418 13666 20428 13819
rect 20494 13666 20504 13819
rect 20610 13666 20620 13819
rect 20686 13666 20696 13819
rect 20802 13666 20812 13819
rect 20878 13666 20888 13819
rect 20994 13666 21004 13819
rect 21070 13666 21080 13819
rect 21186 13666 21196 13819
rect 21262 13666 21272 13819
rect 21378 13666 21388 13819
rect 21454 13666 21464 13819
rect 21570 13666 21580 13819
rect 21636 13666 21816 13819
rect 0 13569 1490 13628
rect 1828 13569 3318 13628
rect 3656 13569 5146 13628
rect 5484 13569 6974 13628
rect 7312 13569 8802 13628
rect 9140 13569 10630 13628
rect 10968 13569 12458 13628
rect 12796 13569 14286 13628
rect 14624 13569 16114 13628
rect 16452 13569 17942 13628
rect 18280 13569 19770 13628
rect 20108 13569 21598 13628
rect 0 13390 1490 13449
rect 1828 13390 3318 13449
rect 3656 13390 5146 13449
rect 5484 13390 6974 13449
rect 7312 13390 8802 13449
rect 9140 13390 10630 13449
rect 10968 13390 12458 13449
rect 12796 13390 14286 13449
rect 14624 13390 16114 13449
rect 16452 13390 17942 13449
rect 18280 13390 19770 13449
rect 20108 13390 21598 13449
rect 22 13165 32 13318
rect 98 13165 108 13318
rect 214 13165 224 13318
rect 290 13165 300 13318
rect 406 13165 416 13318
rect 482 13165 492 13318
rect 598 13165 608 13318
rect 674 13165 684 13318
rect 790 13165 800 13318
rect 866 13165 876 13318
rect 982 13165 992 13318
rect 1058 13165 1068 13318
rect 1174 13165 1184 13318
rect 1250 13165 1260 13318
rect 1366 13165 1376 13318
rect 1442 13165 1452 13318
rect 1488 13105 1708 13352
rect 1850 13165 1860 13318
rect 1926 13165 1936 13318
rect 2042 13165 2052 13318
rect 2118 13165 2128 13318
rect 2234 13165 2244 13318
rect 2310 13165 2320 13318
rect 2426 13165 2436 13318
rect 2502 13165 2512 13318
rect 2618 13165 2628 13318
rect 2694 13165 2704 13318
rect 2810 13165 2820 13318
rect 2886 13165 2896 13318
rect 3002 13165 3012 13318
rect 3078 13165 3088 13318
rect 3194 13165 3204 13318
rect 3270 13165 3280 13318
rect 3316 13105 3536 13352
rect 3678 13165 3688 13318
rect 3754 13165 3764 13318
rect 3870 13165 3880 13318
rect 3946 13165 3956 13318
rect 4062 13165 4072 13318
rect 4138 13165 4148 13318
rect 4254 13165 4264 13318
rect 4330 13165 4340 13318
rect 4446 13165 4456 13318
rect 4522 13165 4532 13318
rect 4638 13165 4648 13318
rect 4714 13165 4724 13318
rect 4830 13165 4840 13318
rect 4906 13165 4916 13318
rect 5022 13165 5032 13318
rect 5098 13165 5108 13318
rect 5144 13105 5364 13352
rect 5506 13165 5516 13318
rect 5582 13165 5592 13318
rect 5698 13165 5708 13318
rect 5774 13165 5784 13318
rect 5890 13165 5900 13318
rect 5966 13165 5976 13318
rect 6082 13165 6092 13318
rect 6158 13165 6168 13318
rect 6274 13165 6284 13318
rect 6350 13165 6360 13318
rect 6466 13165 6476 13318
rect 6542 13165 6552 13318
rect 6658 13165 6668 13318
rect 6734 13165 6744 13318
rect 6850 13165 6860 13318
rect 6926 13165 6936 13318
rect 6972 13105 7192 13352
rect 7334 13165 7344 13318
rect 7410 13165 7420 13318
rect 7526 13165 7536 13318
rect 7602 13165 7612 13318
rect 7718 13165 7728 13318
rect 7794 13165 7804 13318
rect 7910 13165 7920 13318
rect 7986 13165 7996 13318
rect 8102 13165 8112 13318
rect 8178 13165 8188 13318
rect 8294 13165 8304 13318
rect 8370 13165 8380 13318
rect 8486 13165 8496 13318
rect 8562 13165 8572 13318
rect 8678 13165 8688 13318
rect 8754 13165 8764 13318
rect 8800 13105 9020 13352
rect 9162 13165 9172 13318
rect 9238 13165 9248 13318
rect 9354 13165 9364 13318
rect 9430 13165 9440 13318
rect 9546 13165 9556 13318
rect 9622 13165 9632 13318
rect 9738 13165 9748 13318
rect 9814 13165 9824 13318
rect 9930 13165 9940 13318
rect 10006 13165 10016 13318
rect 10122 13165 10132 13318
rect 10198 13165 10208 13318
rect 10314 13165 10324 13318
rect 10390 13165 10400 13318
rect 10506 13165 10516 13318
rect 10582 13165 10592 13318
rect 10628 13105 10848 13352
rect 10990 13165 11000 13318
rect 11066 13165 11076 13318
rect 11182 13165 11192 13318
rect 11258 13165 11268 13318
rect 11374 13165 11384 13318
rect 11450 13165 11460 13318
rect 11566 13165 11576 13318
rect 11642 13165 11652 13318
rect 11758 13165 11768 13318
rect 11834 13165 11844 13318
rect 11950 13165 11960 13318
rect 12026 13165 12036 13318
rect 12142 13165 12152 13318
rect 12218 13165 12228 13318
rect 12334 13165 12344 13318
rect 12410 13165 12420 13318
rect 12456 13105 12676 13352
rect 12818 13165 12828 13318
rect 12894 13165 12904 13318
rect 13010 13165 13020 13318
rect 13086 13165 13096 13318
rect 13202 13165 13212 13318
rect 13278 13165 13288 13318
rect 13394 13165 13404 13318
rect 13470 13165 13480 13318
rect 13586 13165 13596 13318
rect 13662 13165 13672 13318
rect 13778 13165 13788 13318
rect 13854 13165 13864 13318
rect 13970 13165 13980 13318
rect 14046 13165 14056 13318
rect 14162 13165 14172 13318
rect 14238 13165 14248 13318
rect 14284 13105 14504 13352
rect 14646 13165 14656 13318
rect 14722 13165 14732 13318
rect 14838 13165 14848 13318
rect 14914 13165 14924 13318
rect 15030 13165 15040 13318
rect 15106 13165 15116 13318
rect 15222 13165 15232 13318
rect 15298 13165 15308 13318
rect 15414 13165 15424 13318
rect 15490 13165 15500 13318
rect 15606 13165 15616 13318
rect 15682 13165 15692 13318
rect 15798 13165 15808 13318
rect 15874 13165 15884 13318
rect 15990 13165 16000 13318
rect 16066 13165 16076 13318
rect 16112 13105 16332 13352
rect 16474 13165 16484 13318
rect 16550 13165 16560 13318
rect 16666 13165 16676 13318
rect 16742 13165 16752 13318
rect 16858 13165 16868 13318
rect 16934 13165 16944 13318
rect 17050 13165 17060 13318
rect 17126 13165 17136 13318
rect 17242 13165 17252 13318
rect 17318 13165 17328 13318
rect 17434 13165 17444 13318
rect 17510 13165 17520 13318
rect 17626 13165 17636 13318
rect 17702 13165 17712 13318
rect 17818 13165 17828 13318
rect 17894 13165 17904 13318
rect 17940 13105 18160 13352
rect 18302 13165 18312 13318
rect 18378 13165 18388 13318
rect 18494 13165 18504 13318
rect 18570 13165 18580 13318
rect 18686 13165 18696 13318
rect 18762 13165 18772 13318
rect 18878 13165 18888 13318
rect 18954 13165 18964 13318
rect 19070 13165 19080 13318
rect 19146 13165 19156 13318
rect 19262 13165 19272 13318
rect 19338 13165 19348 13318
rect 19454 13165 19464 13318
rect 19530 13165 19540 13318
rect 19646 13165 19656 13318
rect 19722 13165 19732 13318
rect 19768 13105 19988 13352
rect 20130 13165 20140 13318
rect 20206 13165 20216 13318
rect 20322 13165 20332 13318
rect 20398 13165 20408 13318
rect 20514 13165 20524 13318
rect 20590 13165 20600 13318
rect 20706 13165 20716 13318
rect 20782 13165 20792 13318
rect 20898 13165 20908 13318
rect 20974 13165 20984 13318
rect 21090 13165 21100 13318
rect 21166 13165 21176 13318
rect 21282 13165 21292 13318
rect 21358 13165 21368 13318
rect 21474 13165 21484 13318
rect 21550 13165 21560 13318
rect 21596 13105 21816 13352
rect 118 12952 128 13105
rect 194 12952 204 13105
rect 310 12952 320 13105
rect 386 12952 396 13105
rect 502 12952 512 13105
rect 578 12952 588 13105
rect 694 12952 704 13105
rect 770 12952 780 13105
rect 886 12952 896 13105
rect 962 12952 972 13105
rect 1078 12952 1088 13105
rect 1154 12952 1164 13105
rect 1270 12952 1280 13105
rect 1346 12952 1356 13105
rect 1462 12952 1472 13105
rect 1528 12952 1708 13105
rect 1946 12952 1956 13105
rect 2022 12952 2032 13105
rect 2138 12952 2148 13105
rect 2214 12952 2224 13105
rect 2330 12952 2340 13105
rect 2406 12952 2416 13105
rect 2522 12952 2532 13105
rect 2598 12952 2608 13105
rect 2714 12952 2724 13105
rect 2790 12952 2800 13105
rect 2906 12952 2916 13105
rect 2982 12952 2992 13105
rect 3098 12952 3108 13105
rect 3174 12952 3184 13105
rect 3290 12952 3300 13105
rect 3356 12952 3536 13105
rect 3774 12952 3784 13105
rect 3850 12952 3860 13105
rect 3966 12952 3976 13105
rect 4042 12952 4052 13105
rect 4158 12952 4168 13105
rect 4234 12952 4244 13105
rect 4350 12952 4360 13105
rect 4426 12952 4436 13105
rect 4542 12952 4552 13105
rect 4618 12952 4628 13105
rect 4734 12952 4744 13105
rect 4810 12952 4820 13105
rect 4926 12952 4936 13105
rect 5002 12952 5012 13105
rect 5118 12952 5128 13105
rect 5184 12952 5364 13105
rect 5602 12952 5612 13105
rect 5678 12952 5688 13105
rect 5794 12952 5804 13105
rect 5870 12952 5880 13105
rect 5986 12952 5996 13105
rect 6062 12952 6072 13105
rect 6178 12952 6188 13105
rect 6254 12952 6264 13105
rect 6370 12952 6380 13105
rect 6446 12952 6456 13105
rect 6562 12952 6572 13105
rect 6638 12952 6648 13105
rect 6754 12952 6764 13105
rect 6830 12952 6840 13105
rect 6946 12952 6956 13105
rect 7012 12952 7192 13105
rect 7430 12952 7440 13105
rect 7506 12952 7516 13105
rect 7622 12952 7632 13105
rect 7698 12952 7708 13105
rect 7814 12952 7824 13105
rect 7890 12952 7900 13105
rect 8006 12952 8016 13105
rect 8082 12952 8092 13105
rect 8198 12952 8208 13105
rect 8274 12952 8284 13105
rect 8390 12952 8400 13105
rect 8466 12952 8476 13105
rect 8582 12952 8592 13105
rect 8658 12952 8668 13105
rect 8774 12952 8784 13105
rect 8840 12952 9020 13105
rect 9258 12952 9268 13105
rect 9334 12952 9344 13105
rect 9450 12952 9460 13105
rect 9526 12952 9536 13105
rect 9642 12952 9652 13105
rect 9718 12952 9728 13105
rect 9834 12952 9844 13105
rect 9910 12952 9920 13105
rect 10026 12952 10036 13105
rect 10102 12952 10112 13105
rect 10218 12952 10228 13105
rect 10294 12952 10304 13105
rect 10410 12952 10420 13105
rect 10486 12952 10496 13105
rect 10602 12952 10612 13105
rect 10668 12952 10848 13105
rect 11086 12952 11096 13105
rect 11162 12952 11172 13105
rect 11278 12952 11288 13105
rect 11354 12952 11364 13105
rect 11470 12952 11480 13105
rect 11546 12952 11556 13105
rect 11662 12952 11672 13105
rect 11738 12952 11748 13105
rect 11854 12952 11864 13105
rect 11930 12952 11940 13105
rect 12046 12952 12056 13105
rect 12122 12952 12132 13105
rect 12238 12952 12248 13105
rect 12314 12952 12324 13105
rect 12430 12952 12440 13105
rect 12496 12952 12676 13105
rect 12914 12952 12924 13105
rect 12990 12952 13000 13105
rect 13106 12952 13116 13105
rect 13182 12952 13192 13105
rect 13298 12952 13308 13105
rect 13374 12952 13384 13105
rect 13490 12952 13500 13105
rect 13566 12952 13576 13105
rect 13682 12952 13692 13105
rect 13758 12952 13768 13105
rect 13874 12952 13884 13105
rect 13950 12952 13960 13105
rect 14066 12952 14076 13105
rect 14142 12952 14152 13105
rect 14258 12952 14268 13105
rect 14324 12952 14504 13105
rect 14742 12952 14752 13105
rect 14818 12952 14828 13105
rect 14934 12952 14944 13105
rect 15010 12952 15020 13105
rect 15126 12952 15136 13105
rect 15202 12952 15212 13105
rect 15318 12952 15328 13105
rect 15394 12952 15404 13105
rect 15510 12952 15520 13105
rect 15586 12952 15596 13105
rect 15702 12952 15712 13105
rect 15778 12952 15788 13105
rect 15894 12952 15904 13105
rect 15970 12952 15980 13105
rect 16086 12952 16096 13105
rect 16152 12952 16332 13105
rect 16570 12952 16580 13105
rect 16646 12952 16656 13105
rect 16762 12952 16772 13105
rect 16838 12952 16848 13105
rect 16954 12952 16964 13105
rect 17030 12952 17040 13105
rect 17146 12952 17156 13105
rect 17222 12952 17232 13105
rect 17338 12952 17348 13105
rect 17414 12952 17424 13105
rect 17530 12952 17540 13105
rect 17606 12952 17616 13105
rect 17722 12952 17732 13105
rect 17798 12952 17808 13105
rect 17914 12952 17924 13105
rect 17980 12952 18160 13105
rect 18398 12952 18408 13105
rect 18474 12952 18484 13105
rect 18590 12952 18600 13105
rect 18666 12952 18676 13105
rect 18782 12952 18792 13105
rect 18858 12952 18868 13105
rect 18974 12952 18984 13105
rect 19050 12952 19060 13105
rect 19166 12952 19176 13105
rect 19242 12952 19252 13105
rect 19358 12952 19368 13105
rect 19434 12952 19444 13105
rect 19550 12952 19560 13105
rect 19626 12952 19636 13105
rect 19742 12952 19752 13105
rect 19808 12952 19988 13105
rect 20226 12952 20236 13105
rect 20302 12952 20312 13105
rect 20418 12952 20428 13105
rect 20494 12952 20504 13105
rect 20610 12952 20620 13105
rect 20686 12952 20696 13105
rect 20802 12952 20812 13105
rect 20878 12952 20888 13105
rect 20994 12952 21004 13105
rect 21070 12952 21080 13105
rect 21186 12952 21196 13105
rect 21262 12952 21272 13105
rect 21378 12952 21388 13105
rect 21454 12952 21464 13105
rect 21570 12952 21580 13105
rect 21636 12952 21816 13105
rect 0 12855 1490 12914
rect 1828 12855 3318 12914
rect 3656 12855 5146 12914
rect 5484 12855 6974 12914
rect 7312 12855 8802 12914
rect 9140 12855 10630 12914
rect 10968 12855 12458 12914
rect 12796 12855 14286 12914
rect 14624 12855 16114 12914
rect 16452 12855 17942 12914
rect 18280 12855 19770 12914
rect 20108 12855 21598 12914
rect 0 12676 1490 12735
rect 1828 12676 3318 12735
rect 3656 12676 5146 12735
rect 5484 12676 6974 12735
rect 7312 12676 8802 12735
rect 9140 12676 10630 12735
rect 10968 12676 12458 12735
rect 12796 12676 14286 12735
rect 14624 12676 16114 12735
rect 16452 12676 17942 12735
rect 18280 12676 19770 12735
rect 20108 12676 21598 12735
rect 22 12451 32 12604
rect 98 12451 108 12604
rect 214 12451 224 12604
rect 290 12451 300 12604
rect 406 12451 416 12604
rect 482 12451 492 12604
rect 598 12451 608 12604
rect 674 12451 684 12604
rect 790 12451 800 12604
rect 866 12451 876 12604
rect 982 12451 992 12604
rect 1058 12451 1068 12604
rect 1174 12451 1184 12604
rect 1250 12451 1260 12604
rect 1366 12451 1376 12604
rect 1442 12451 1452 12604
rect 1488 12391 1708 12638
rect 1850 12451 1860 12604
rect 1926 12451 1936 12604
rect 2042 12451 2052 12604
rect 2118 12451 2128 12604
rect 2234 12451 2244 12604
rect 2310 12451 2320 12604
rect 2426 12451 2436 12604
rect 2502 12451 2512 12604
rect 2618 12451 2628 12604
rect 2694 12451 2704 12604
rect 2810 12451 2820 12604
rect 2886 12451 2896 12604
rect 3002 12451 3012 12604
rect 3078 12451 3088 12604
rect 3194 12451 3204 12604
rect 3270 12451 3280 12604
rect 3316 12391 3536 12638
rect 3678 12451 3688 12604
rect 3754 12451 3764 12604
rect 3870 12451 3880 12604
rect 3946 12451 3956 12604
rect 4062 12451 4072 12604
rect 4138 12451 4148 12604
rect 4254 12451 4264 12604
rect 4330 12451 4340 12604
rect 4446 12451 4456 12604
rect 4522 12451 4532 12604
rect 4638 12451 4648 12604
rect 4714 12451 4724 12604
rect 4830 12451 4840 12604
rect 4906 12451 4916 12604
rect 5022 12451 5032 12604
rect 5098 12451 5108 12604
rect 5144 12391 5364 12638
rect 5506 12451 5516 12604
rect 5582 12451 5592 12604
rect 5698 12451 5708 12604
rect 5774 12451 5784 12604
rect 5890 12451 5900 12604
rect 5966 12451 5976 12604
rect 6082 12451 6092 12604
rect 6158 12451 6168 12604
rect 6274 12451 6284 12604
rect 6350 12451 6360 12604
rect 6466 12451 6476 12604
rect 6542 12451 6552 12604
rect 6658 12451 6668 12604
rect 6734 12451 6744 12604
rect 6850 12451 6860 12604
rect 6926 12451 6936 12604
rect 6972 12391 7192 12638
rect 7334 12451 7344 12604
rect 7410 12451 7420 12604
rect 7526 12451 7536 12604
rect 7602 12451 7612 12604
rect 7718 12451 7728 12604
rect 7794 12451 7804 12604
rect 7910 12451 7920 12604
rect 7986 12451 7996 12604
rect 8102 12451 8112 12604
rect 8178 12451 8188 12604
rect 8294 12451 8304 12604
rect 8370 12451 8380 12604
rect 8486 12451 8496 12604
rect 8562 12451 8572 12604
rect 8678 12451 8688 12604
rect 8754 12451 8764 12604
rect 8800 12391 9020 12638
rect 9162 12451 9172 12604
rect 9238 12451 9248 12604
rect 9354 12451 9364 12604
rect 9430 12451 9440 12604
rect 9546 12451 9556 12604
rect 9622 12451 9632 12604
rect 9738 12451 9748 12604
rect 9814 12451 9824 12604
rect 9930 12451 9940 12604
rect 10006 12451 10016 12604
rect 10122 12451 10132 12604
rect 10198 12451 10208 12604
rect 10314 12451 10324 12604
rect 10390 12451 10400 12604
rect 10506 12451 10516 12604
rect 10582 12451 10592 12604
rect 10628 12391 10848 12638
rect 10990 12451 11000 12604
rect 11066 12451 11076 12604
rect 11182 12451 11192 12604
rect 11258 12451 11268 12604
rect 11374 12451 11384 12604
rect 11450 12451 11460 12604
rect 11566 12451 11576 12604
rect 11642 12451 11652 12604
rect 11758 12451 11768 12604
rect 11834 12451 11844 12604
rect 11950 12451 11960 12604
rect 12026 12451 12036 12604
rect 12142 12451 12152 12604
rect 12218 12451 12228 12604
rect 12334 12451 12344 12604
rect 12410 12451 12420 12604
rect 12456 12391 12676 12638
rect 12818 12451 12828 12604
rect 12894 12451 12904 12604
rect 13010 12451 13020 12604
rect 13086 12451 13096 12604
rect 13202 12451 13212 12604
rect 13278 12451 13288 12604
rect 13394 12451 13404 12604
rect 13470 12451 13480 12604
rect 13586 12451 13596 12604
rect 13662 12451 13672 12604
rect 13778 12451 13788 12604
rect 13854 12451 13864 12604
rect 13970 12451 13980 12604
rect 14046 12451 14056 12604
rect 14162 12451 14172 12604
rect 14238 12451 14248 12604
rect 14284 12391 14504 12638
rect 14646 12451 14656 12604
rect 14722 12451 14732 12604
rect 14838 12451 14848 12604
rect 14914 12451 14924 12604
rect 15030 12451 15040 12604
rect 15106 12451 15116 12604
rect 15222 12451 15232 12604
rect 15298 12451 15308 12604
rect 15414 12451 15424 12604
rect 15490 12451 15500 12604
rect 15606 12451 15616 12604
rect 15682 12451 15692 12604
rect 15798 12451 15808 12604
rect 15874 12451 15884 12604
rect 15990 12451 16000 12604
rect 16066 12451 16076 12604
rect 16112 12391 16332 12638
rect 16474 12451 16484 12604
rect 16550 12451 16560 12604
rect 16666 12451 16676 12604
rect 16742 12451 16752 12604
rect 16858 12451 16868 12604
rect 16934 12451 16944 12604
rect 17050 12451 17060 12604
rect 17126 12451 17136 12604
rect 17242 12451 17252 12604
rect 17318 12451 17328 12604
rect 17434 12451 17444 12604
rect 17510 12451 17520 12604
rect 17626 12451 17636 12604
rect 17702 12451 17712 12604
rect 17818 12451 17828 12604
rect 17894 12451 17904 12604
rect 17940 12391 18160 12638
rect 18302 12451 18312 12604
rect 18378 12451 18388 12604
rect 18494 12451 18504 12604
rect 18570 12451 18580 12604
rect 18686 12451 18696 12604
rect 18762 12451 18772 12604
rect 18878 12451 18888 12604
rect 18954 12451 18964 12604
rect 19070 12451 19080 12604
rect 19146 12451 19156 12604
rect 19262 12451 19272 12604
rect 19338 12451 19348 12604
rect 19454 12451 19464 12604
rect 19530 12451 19540 12604
rect 19646 12451 19656 12604
rect 19722 12451 19732 12604
rect 19768 12391 19988 12638
rect 20130 12451 20140 12604
rect 20206 12451 20216 12604
rect 20322 12451 20332 12604
rect 20398 12451 20408 12604
rect 20514 12451 20524 12604
rect 20590 12451 20600 12604
rect 20706 12451 20716 12604
rect 20782 12451 20792 12604
rect 20898 12451 20908 12604
rect 20974 12451 20984 12604
rect 21090 12451 21100 12604
rect 21166 12451 21176 12604
rect 21282 12451 21292 12604
rect 21358 12451 21368 12604
rect 21474 12451 21484 12604
rect 21550 12451 21560 12604
rect 21596 12391 21816 12638
rect 118 12238 128 12391
rect 194 12238 204 12391
rect 310 12238 320 12391
rect 386 12238 396 12391
rect 502 12238 512 12391
rect 578 12238 588 12391
rect 694 12238 704 12391
rect 770 12238 780 12391
rect 886 12238 896 12391
rect 962 12238 972 12391
rect 1078 12238 1088 12391
rect 1154 12238 1164 12391
rect 1270 12238 1280 12391
rect 1346 12238 1356 12391
rect 1462 12238 1472 12391
rect 1528 12238 1708 12391
rect 1946 12238 1956 12391
rect 2022 12238 2032 12391
rect 2138 12238 2148 12391
rect 2214 12238 2224 12391
rect 2330 12238 2340 12391
rect 2406 12238 2416 12391
rect 2522 12238 2532 12391
rect 2598 12238 2608 12391
rect 2714 12238 2724 12391
rect 2790 12238 2800 12391
rect 2906 12238 2916 12391
rect 2982 12238 2992 12391
rect 3098 12238 3108 12391
rect 3174 12238 3184 12391
rect 3290 12238 3300 12391
rect 3356 12238 3536 12391
rect 3774 12238 3784 12391
rect 3850 12238 3860 12391
rect 3966 12238 3976 12391
rect 4042 12238 4052 12391
rect 4158 12238 4168 12391
rect 4234 12238 4244 12391
rect 4350 12238 4360 12391
rect 4426 12238 4436 12391
rect 4542 12238 4552 12391
rect 4618 12238 4628 12391
rect 4734 12238 4744 12391
rect 4810 12238 4820 12391
rect 4926 12238 4936 12391
rect 5002 12238 5012 12391
rect 5118 12238 5128 12391
rect 5184 12238 5364 12391
rect 5602 12238 5612 12391
rect 5678 12238 5688 12391
rect 5794 12238 5804 12391
rect 5870 12238 5880 12391
rect 5986 12238 5996 12391
rect 6062 12238 6072 12391
rect 6178 12238 6188 12391
rect 6254 12238 6264 12391
rect 6370 12238 6380 12391
rect 6446 12238 6456 12391
rect 6562 12238 6572 12391
rect 6638 12238 6648 12391
rect 6754 12238 6764 12391
rect 6830 12238 6840 12391
rect 6946 12238 6956 12391
rect 7012 12238 7192 12391
rect 7430 12238 7440 12391
rect 7506 12238 7516 12391
rect 7622 12238 7632 12391
rect 7698 12238 7708 12391
rect 7814 12238 7824 12391
rect 7890 12238 7900 12391
rect 8006 12238 8016 12391
rect 8082 12238 8092 12391
rect 8198 12238 8208 12391
rect 8274 12238 8284 12391
rect 8390 12238 8400 12391
rect 8466 12238 8476 12391
rect 8582 12238 8592 12391
rect 8658 12238 8668 12391
rect 8774 12238 8784 12391
rect 8840 12238 9020 12391
rect 9258 12238 9268 12391
rect 9334 12238 9344 12391
rect 9450 12238 9460 12391
rect 9526 12238 9536 12391
rect 9642 12238 9652 12391
rect 9718 12238 9728 12391
rect 9834 12238 9844 12391
rect 9910 12238 9920 12391
rect 10026 12238 10036 12391
rect 10102 12238 10112 12391
rect 10218 12238 10228 12391
rect 10294 12238 10304 12391
rect 10410 12238 10420 12391
rect 10486 12238 10496 12391
rect 10602 12238 10612 12391
rect 10668 12238 10848 12391
rect 11086 12238 11096 12391
rect 11162 12238 11172 12391
rect 11278 12238 11288 12391
rect 11354 12238 11364 12391
rect 11470 12238 11480 12391
rect 11546 12238 11556 12391
rect 11662 12238 11672 12391
rect 11738 12238 11748 12391
rect 11854 12238 11864 12391
rect 11930 12238 11940 12391
rect 12046 12238 12056 12391
rect 12122 12238 12132 12391
rect 12238 12238 12248 12391
rect 12314 12238 12324 12391
rect 12430 12238 12440 12391
rect 12496 12238 12676 12391
rect 12914 12238 12924 12391
rect 12990 12238 13000 12391
rect 13106 12238 13116 12391
rect 13182 12238 13192 12391
rect 13298 12238 13308 12391
rect 13374 12238 13384 12391
rect 13490 12238 13500 12391
rect 13566 12238 13576 12391
rect 13682 12238 13692 12391
rect 13758 12238 13768 12391
rect 13874 12238 13884 12391
rect 13950 12238 13960 12391
rect 14066 12238 14076 12391
rect 14142 12238 14152 12391
rect 14258 12238 14268 12391
rect 14324 12238 14504 12391
rect 14742 12238 14752 12391
rect 14818 12238 14828 12391
rect 14934 12238 14944 12391
rect 15010 12238 15020 12391
rect 15126 12238 15136 12391
rect 15202 12238 15212 12391
rect 15318 12238 15328 12391
rect 15394 12238 15404 12391
rect 15510 12238 15520 12391
rect 15586 12238 15596 12391
rect 15702 12238 15712 12391
rect 15778 12238 15788 12391
rect 15894 12238 15904 12391
rect 15970 12238 15980 12391
rect 16086 12238 16096 12391
rect 16152 12238 16332 12391
rect 16570 12238 16580 12391
rect 16646 12238 16656 12391
rect 16762 12238 16772 12391
rect 16838 12238 16848 12391
rect 16954 12238 16964 12391
rect 17030 12238 17040 12391
rect 17146 12238 17156 12391
rect 17222 12238 17232 12391
rect 17338 12238 17348 12391
rect 17414 12238 17424 12391
rect 17530 12238 17540 12391
rect 17606 12238 17616 12391
rect 17722 12238 17732 12391
rect 17798 12238 17808 12391
rect 17914 12238 17924 12391
rect 17980 12238 18160 12391
rect 18398 12238 18408 12391
rect 18474 12238 18484 12391
rect 18590 12238 18600 12391
rect 18666 12238 18676 12391
rect 18782 12238 18792 12391
rect 18858 12238 18868 12391
rect 18974 12238 18984 12391
rect 19050 12238 19060 12391
rect 19166 12238 19176 12391
rect 19242 12238 19252 12391
rect 19358 12238 19368 12391
rect 19434 12238 19444 12391
rect 19550 12238 19560 12391
rect 19626 12238 19636 12391
rect 19742 12238 19752 12391
rect 19808 12238 19988 12391
rect 20226 12238 20236 12391
rect 20302 12238 20312 12391
rect 20418 12238 20428 12391
rect 20494 12238 20504 12391
rect 20610 12238 20620 12391
rect 20686 12238 20696 12391
rect 20802 12238 20812 12391
rect 20878 12238 20888 12391
rect 20994 12238 21004 12391
rect 21070 12238 21080 12391
rect 21186 12238 21196 12391
rect 21262 12238 21272 12391
rect 21378 12238 21388 12391
rect 21454 12238 21464 12391
rect 21570 12238 21580 12391
rect 21636 12238 21816 12391
rect 0 12141 1490 12200
rect 1828 12141 3318 12200
rect 3656 12141 5146 12200
rect 5484 12141 6974 12200
rect 7312 12141 8802 12200
rect 9140 12141 10630 12200
rect 10968 12141 12458 12200
rect 12796 12141 14286 12200
rect 14624 12141 16114 12200
rect 16452 12141 17942 12200
rect 18280 12141 19770 12200
rect 20108 12141 21598 12200
rect 0 11962 1490 12021
rect 1828 11962 3318 12021
rect 3656 11962 5146 12021
rect 5484 11962 6974 12021
rect 7312 11962 8802 12021
rect 9140 11962 10630 12021
rect 10968 11962 12458 12021
rect 12796 11962 14286 12021
rect 14624 11962 16114 12021
rect 16452 11962 17942 12021
rect 18280 11962 19770 12021
rect 20108 11962 21598 12021
rect 22 11737 32 11890
rect 98 11737 108 11890
rect 214 11737 224 11890
rect 290 11737 300 11890
rect 406 11737 416 11890
rect 482 11737 492 11890
rect 598 11737 608 11890
rect 674 11737 684 11890
rect 790 11737 800 11890
rect 866 11737 876 11890
rect 982 11737 992 11890
rect 1058 11737 1068 11890
rect 1174 11737 1184 11890
rect 1250 11737 1260 11890
rect 1366 11737 1376 11890
rect 1442 11737 1452 11890
rect 1488 11677 1708 11924
rect 1850 11737 1860 11890
rect 1926 11737 1936 11890
rect 2042 11737 2052 11890
rect 2118 11737 2128 11890
rect 2234 11737 2244 11890
rect 2310 11737 2320 11890
rect 2426 11737 2436 11890
rect 2502 11737 2512 11890
rect 2618 11737 2628 11890
rect 2694 11737 2704 11890
rect 2810 11737 2820 11890
rect 2886 11737 2896 11890
rect 3002 11737 3012 11890
rect 3078 11737 3088 11890
rect 3194 11737 3204 11890
rect 3270 11737 3280 11890
rect 3316 11677 3536 11924
rect 3678 11737 3688 11890
rect 3754 11737 3764 11890
rect 3870 11737 3880 11890
rect 3946 11737 3956 11890
rect 4062 11737 4072 11890
rect 4138 11737 4148 11890
rect 4254 11737 4264 11890
rect 4330 11737 4340 11890
rect 4446 11737 4456 11890
rect 4522 11737 4532 11890
rect 4638 11737 4648 11890
rect 4714 11737 4724 11890
rect 4830 11737 4840 11890
rect 4906 11737 4916 11890
rect 5022 11737 5032 11890
rect 5098 11737 5108 11890
rect 5144 11677 5364 11924
rect 5506 11737 5516 11890
rect 5582 11737 5592 11890
rect 5698 11737 5708 11890
rect 5774 11737 5784 11890
rect 5890 11737 5900 11890
rect 5966 11737 5976 11890
rect 6082 11737 6092 11890
rect 6158 11737 6168 11890
rect 6274 11737 6284 11890
rect 6350 11737 6360 11890
rect 6466 11737 6476 11890
rect 6542 11737 6552 11890
rect 6658 11737 6668 11890
rect 6734 11737 6744 11890
rect 6850 11737 6860 11890
rect 6926 11737 6936 11890
rect 6972 11677 7192 11924
rect 7334 11737 7344 11890
rect 7410 11737 7420 11890
rect 7526 11737 7536 11890
rect 7602 11737 7612 11890
rect 7718 11737 7728 11890
rect 7794 11737 7804 11890
rect 7910 11737 7920 11890
rect 7986 11737 7996 11890
rect 8102 11737 8112 11890
rect 8178 11737 8188 11890
rect 8294 11737 8304 11890
rect 8370 11737 8380 11890
rect 8486 11737 8496 11890
rect 8562 11737 8572 11890
rect 8678 11737 8688 11890
rect 8754 11737 8764 11890
rect 8800 11677 9020 11924
rect 9162 11737 9172 11890
rect 9238 11737 9248 11890
rect 9354 11737 9364 11890
rect 9430 11737 9440 11890
rect 9546 11737 9556 11890
rect 9622 11737 9632 11890
rect 9738 11737 9748 11890
rect 9814 11737 9824 11890
rect 9930 11737 9940 11890
rect 10006 11737 10016 11890
rect 10122 11737 10132 11890
rect 10198 11737 10208 11890
rect 10314 11737 10324 11890
rect 10390 11737 10400 11890
rect 10506 11737 10516 11890
rect 10582 11737 10592 11890
rect 10628 11677 10848 11924
rect 10990 11737 11000 11890
rect 11066 11737 11076 11890
rect 11182 11737 11192 11890
rect 11258 11737 11268 11890
rect 11374 11737 11384 11890
rect 11450 11737 11460 11890
rect 11566 11737 11576 11890
rect 11642 11737 11652 11890
rect 11758 11737 11768 11890
rect 11834 11737 11844 11890
rect 11950 11737 11960 11890
rect 12026 11737 12036 11890
rect 12142 11737 12152 11890
rect 12218 11737 12228 11890
rect 12334 11737 12344 11890
rect 12410 11737 12420 11890
rect 12456 11677 12676 11924
rect 12818 11737 12828 11890
rect 12894 11737 12904 11890
rect 13010 11737 13020 11890
rect 13086 11737 13096 11890
rect 13202 11737 13212 11890
rect 13278 11737 13288 11890
rect 13394 11737 13404 11890
rect 13470 11737 13480 11890
rect 13586 11737 13596 11890
rect 13662 11737 13672 11890
rect 13778 11737 13788 11890
rect 13854 11737 13864 11890
rect 13970 11737 13980 11890
rect 14046 11737 14056 11890
rect 14162 11737 14172 11890
rect 14238 11737 14248 11890
rect 14284 11677 14504 11924
rect 14646 11737 14656 11890
rect 14722 11737 14732 11890
rect 14838 11737 14848 11890
rect 14914 11737 14924 11890
rect 15030 11737 15040 11890
rect 15106 11737 15116 11890
rect 15222 11737 15232 11890
rect 15298 11737 15308 11890
rect 15414 11737 15424 11890
rect 15490 11737 15500 11890
rect 15606 11737 15616 11890
rect 15682 11737 15692 11890
rect 15798 11737 15808 11890
rect 15874 11737 15884 11890
rect 15990 11737 16000 11890
rect 16066 11737 16076 11890
rect 16112 11677 16332 11924
rect 16474 11737 16484 11890
rect 16550 11737 16560 11890
rect 16666 11737 16676 11890
rect 16742 11737 16752 11890
rect 16858 11737 16868 11890
rect 16934 11737 16944 11890
rect 17050 11737 17060 11890
rect 17126 11737 17136 11890
rect 17242 11737 17252 11890
rect 17318 11737 17328 11890
rect 17434 11737 17444 11890
rect 17510 11737 17520 11890
rect 17626 11737 17636 11890
rect 17702 11737 17712 11890
rect 17818 11737 17828 11890
rect 17894 11737 17904 11890
rect 17940 11677 18160 11924
rect 18302 11737 18312 11890
rect 18378 11737 18388 11890
rect 18494 11737 18504 11890
rect 18570 11737 18580 11890
rect 18686 11737 18696 11890
rect 18762 11737 18772 11890
rect 18878 11737 18888 11890
rect 18954 11737 18964 11890
rect 19070 11737 19080 11890
rect 19146 11737 19156 11890
rect 19262 11737 19272 11890
rect 19338 11737 19348 11890
rect 19454 11737 19464 11890
rect 19530 11737 19540 11890
rect 19646 11737 19656 11890
rect 19722 11737 19732 11890
rect 19768 11677 19988 11924
rect 20130 11737 20140 11890
rect 20206 11737 20216 11890
rect 20322 11737 20332 11890
rect 20398 11737 20408 11890
rect 20514 11737 20524 11890
rect 20590 11737 20600 11890
rect 20706 11737 20716 11890
rect 20782 11737 20792 11890
rect 20898 11737 20908 11890
rect 20974 11737 20984 11890
rect 21090 11737 21100 11890
rect 21166 11737 21176 11890
rect 21282 11737 21292 11890
rect 21358 11737 21368 11890
rect 21474 11737 21484 11890
rect 21550 11737 21560 11890
rect 21596 11677 21816 11924
rect 118 11524 128 11677
rect 194 11524 204 11677
rect 310 11524 320 11677
rect 386 11524 396 11677
rect 502 11524 512 11677
rect 578 11524 588 11677
rect 694 11524 704 11677
rect 770 11524 780 11677
rect 886 11524 896 11677
rect 962 11524 972 11677
rect 1078 11524 1088 11677
rect 1154 11524 1164 11677
rect 1270 11524 1280 11677
rect 1346 11524 1356 11677
rect 1462 11524 1472 11677
rect 1528 11524 1708 11677
rect 1946 11524 1956 11677
rect 2022 11524 2032 11677
rect 2138 11524 2148 11677
rect 2214 11524 2224 11677
rect 2330 11524 2340 11677
rect 2406 11524 2416 11677
rect 2522 11524 2532 11677
rect 2598 11524 2608 11677
rect 2714 11524 2724 11677
rect 2790 11524 2800 11677
rect 2906 11524 2916 11677
rect 2982 11524 2992 11677
rect 3098 11524 3108 11677
rect 3174 11524 3184 11677
rect 3290 11524 3300 11677
rect 3356 11524 3536 11677
rect 3774 11524 3784 11677
rect 3850 11524 3860 11677
rect 3966 11524 3976 11677
rect 4042 11524 4052 11677
rect 4158 11524 4168 11677
rect 4234 11524 4244 11677
rect 4350 11524 4360 11677
rect 4426 11524 4436 11677
rect 4542 11524 4552 11677
rect 4618 11524 4628 11677
rect 4734 11524 4744 11677
rect 4810 11524 4820 11677
rect 4926 11524 4936 11677
rect 5002 11524 5012 11677
rect 5118 11524 5128 11677
rect 5184 11524 5364 11677
rect 5602 11524 5612 11677
rect 5678 11524 5688 11677
rect 5794 11524 5804 11677
rect 5870 11524 5880 11677
rect 5986 11524 5996 11677
rect 6062 11524 6072 11677
rect 6178 11524 6188 11677
rect 6254 11524 6264 11677
rect 6370 11524 6380 11677
rect 6446 11524 6456 11677
rect 6562 11524 6572 11677
rect 6638 11524 6648 11677
rect 6754 11524 6764 11677
rect 6830 11524 6840 11677
rect 6946 11524 6956 11677
rect 7012 11524 7192 11677
rect 7430 11524 7440 11677
rect 7506 11524 7516 11677
rect 7622 11524 7632 11677
rect 7698 11524 7708 11677
rect 7814 11524 7824 11677
rect 7890 11524 7900 11677
rect 8006 11524 8016 11677
rect 8082 11524 8092 11677
rect 8198 11524 8208 11677
rect 8274 11524 8284 11677
rect 8390 11524 8400 11677
rect 8466 11524 8476 11677
rect 8582 11524 8592 11677
rect 8658 11524 8668 11677
rect 8774 11524 8784 11677
rect 8840 11524 9020 11677
rect 9258 11524 9268 11677
rect 9334 11524 9344 11677
rect 9450 11524 9460 11677
rect 9526 11524 9536 11677
rect 9642 11524 9652 11677
rect 9718 11524 9728 11677
rect 9834 11524 9844 11677
rect 9910 11524 9920 11677
rect 10026 11524 10036 11677
rect 10102 11524 10112 11677
rect 10218 11524 10228 11677
rect 10294 11524 10304 11677
rect 10410 11524 10420 11677
rect 10486 11524 10496 11677
rect 10602 11524 10612 11677
rect 10668 11524 10848 11677
rect 11086 11524 11096 11677
rect 11162 11524 11172 11677
rect 11278 11524 11288 11677
rect 11354 11524 11364 11677
rect 11470 11524 11480 11677
rect 11546 11524 11556 11677
rect 11662 11524 11672 11677
rect 11738 11524 11748 11677
rect 11854 11524 11864 11677
rect 11930 11524 11940 11677
rect 12046 11524 12056 11677
rect 12122 11524 12132 11677
rect 12238 11524 12248 11677
rect 12314 11524 12324 11677
rect 12430 11524 12440 11677
rect 12496 11524 12676 11677
rect 12914 11524 12924 11677
rect 12990 11524 13000 11677
rect 13106 11524 13116 11677
rect 13182 11524 13192 11677
rect 13298 11524 13308 11677
rect 13374 11524 13384 11677
rect 13490 11524 13500 11677
rect 13566 11524 13576 11677
rect 13682 11524 13692 11677
rect 13758 11524 13768 11677
rect 13874 11524 13884 11677
rect 13950 11524 13960 11677
rect 14066 11524 14076 11677
rect 14142 11524 14152 11677
rect 14258 11524 14268 11677
rect 14324 11524 14504 11677
rect 14742 11524 14752 11677
rect 14818 11524 14828 11677
rect 14934 11524 14944 11677
rect 15010 11524 15020 11677
rect 15126 11524 15136 11677
rect 15202 11524 15212 11677
rect 15318 11524 15328 11677
rect 15394 11524 15404 11677
rect 15510 11524 15520 11677
rect 15586 11524 15596 11677
rect 15702 11524 15712 11677
rect 15778 11524 15788 11677
rect 15894 11524 15904 11677
rect 15970 11524 15980 11677
rect 16086 11524 16096 11677
rect 16152 11524 16332 11677
rect 16570 11524 16580 11677
rect 16646 11524 16656 11677
rect 16762 11524 16772 11677
rect 16838 11524 16848 11677
rect 16954 11524 16964 11677
rect 17030 11524 17040 11677
rect 17146 11524 17156 11677
rect 17222 11524 17232 11677
rect 17338 11524 17348 11677
rect 17414 11524 17424 11677
rect 17530 11524 17540 11677
rect 17606 11524 17616 11677
rect 17722 11524 17732 11677
rect 17798 11524 17808 11677
rect 17914 11524 17924 11677
rect 17980 11524 18160 11677
rect 18398 11524 18408 11677
rect 18474 11524 18484 11677
rect 18590 11524 18600 11677
rect 18666 11524 18676 11677
rect 18782 11524 18792 11677
rect 18858 11524 18868 11677
rect 18974 11524 18984 11677
rect 19050 11524 19060 11677
rect 19166 11524 19176 11677
rect 19242 11524 19252 11677
rect 19358 11524 19368 11677
rect 19434 11524 19444 11677
rect 19550 11524 19560 11677
rect 19626 11524 19636 11677
rect 19742 11524 19752 11677
rect 19808 11524 19988 11677
rect 20226 11524 20236 11677
rect 20302 11524 20312 11677
rect 20418 11524 20428 11677
rect 20494 11524 20504 11677
rect 20610 11524 20620 11677
rect 20686 11524 20696 11677
rect 20802 11524 20812 11677
rect 20878 11524 20888 11677
rect 20994 11524 21004 11677
rect 21070 11524 21080 11677
rect 21186 11524 21196 11677
rect 21262 11524 21272 11677
rect 21378 11524 21388 11677
rect 21454 11524 21464 11677
rect 21570 11524 21580 11677
rect 21636 11524 21816 11677
rect 0 11427 1490 11486
rect 1828 11427 3318 11486
rect 3656 11427 5146 11486
rect 5484 11427 6974 11486
rect 7312 11427 8802 11486
rect 9140 11427 10630 11486
rect 10968 11427 12458 11486
rect 12796 11427 14286 11486
rect 14624 11427 16114 11486
rect 16452 11427 17942 11486
rect 18280 11427 19770 11486
rect 20108 11427 21598 11486
rect 0 11248 1490 11307
rect 1828 11248 3318 11307
rect 3656 11248 5146 11307
rect 5484 11248 6974 11307
rect 7312 11248 8802 11307
rect 9140 11248 10630 11307
rect 10968 11248 12458 11307
rect 12796 11248 14286 11307
rect 14624 11248 16114 11307
rect 16452 11248 17942 11307
rect 18280 11248 19770 11307
rect 20108 11248 21598 11307
rect 22 11023 32 11176
rect 98 11023 108 11176
rect 214 11023 224 11176
rect 290 11023 300 11176
rect 406 11023 416 11176
rect 482 11023 492 11176
rect 598 11023 608 11176
rect 674 11023 684 11176
rect 790 11023 800 11176
rect 866 11023 876 11176
rect 982 11023 992 11176
rect 1058 11023 1068 11176
rect 1174 11023 1184 11176
rect 1250 11023 1260 11176
rect 1366 11023 1376 11176
rect 1442 11023 1452 11176
rect 1488 10963 1708 11210
rect 1850 11023 1860 11176
rect 1926 11023 1936 11176
rect 2042 11023 2052 11176
rect 2118 11023 2128 11176
rect 2234 11023 2244 11176
rect 2310 11023 2320 11176
rect 2426 11023 2436 11176
rect 2502 11023 2512 11176
rect 2618 11023 2628 11176
rect 2694 11023 2704 11176
rect 2810 11023 2820 11176
rect 2886 11023 2896 11176
rect 3002 11023 3012 11176
rect 3078 11023 3088 11176
rect 3194 11023 3204 11176
rect 3270 11023 3280 11176
rect 3316 10963 3536 11210
rect 3678 11023 3688 11176
rect 3754 11023 3764 11176
rect 3870 11023 3880 11176
rect 3946 11023 3956 11176
rect 4062 11023 4072 11176
rect 4138 11023 4148 11176
rect 4254 11023 4264 11176
rect 4330 11023 4340 11176
rect 4446 11023 4456 11176
rect 4522 11023 4532 11176
rect 4638 11023 4648 11176
rect 4714 11023 4724 11176
rect 4830 11023 4840 11176
rect 4906 11023 4916 11176
rect 5022 11023 5032 11176
rect 5098 11023 5108 11176
rect 5144 10963 5364 11210
rect 5506 11023 5516 11176
rect 5582 11023 5592 11176
rect 5698 11023 5708 11176
rect 5774 11023 5784 11176
rect 5890 11023 5900 11176
rect 5966 11023 5976 11176
rect 6082 11023 6092 11176
rect 6158 11023 6168 11176
rect 6274 11023 6284 11176
rect 6350 11023 6360 11176
rect 6466 11023 6476 11176
rect 6542 11023 6552 11176
rect 6658 11023 6668 11176
rect 6734 11023 6744 11176
rect 6850 11023 6860 11176
rect 6926 11023 6936 11176
rect 6972 10963 7192 11210
rect 7334 11023 7344 11176
rect 7410 11023 7420 11176
rect 7526 11023 7536 11176
rect 7602 11023 7612 11176
rect 7718 11023 7728 11176
rect 7794 11023 7804 11176
rect 7910 11023 7920 11176
rect 7986 11023 7996 11176
rect 8102 11023 8112 11176
rect 8178 11023 8188 11176
rect 8294 11023 8304 11176
rect 8370 11023 8380 11176
rect 8486 11023 8496 11176
rect 8562 11023 8572 11176
rect 8678 11023 8688 11176
rect 8754 11023 8764 11176
rect 8800 10963 9020 11210
rect 9162 11023 9172 11176
rect 9238 11023 9248 11176
rect 9354 11023 9364 11176
rect 9430 11023 9440 11176
rect 9546 11023 9556 11176
rect 9622 11023 9632 11176
rect 9738 11023 9748 11176
rect 9814 11023 9824 11176
rect 9930 11023 9940 11176
rect 10006 11023 10016 11176
rect 10122 11023 10132 11176
rect 10198 11023 10208 11176
rect 10314 11023 10324 11176
rect 10390 11023 10400 11176
rect 10506 11023 10516 11176
rect 10582 11023 10592 11176
rect 10628 10963 10848 11210
rect 10990 11023 11000 11176
rect 11066 11023 11076 11176
rect 11182 11023 11192 11176
rect 11258 11023 11268 11176
rect 11374 11023 11384 11176
rect 11450 11023 11460 11176
rect 11566 11023 11576 11176
rect 11642 11023 11652 11176
rect 11758 11023 11768 11176
rect 11834 11023 11844 11176
rect 11950 11023 11960 11176
rect 12026 11023 12036 11176
rect 12142 11023 12152 11176
rect 12218 11023 12228 11176
rect 12334 11023 12344 11176
rect 12410 11023 12420 11176
rect 12456 10963 12676 11210
rect 12818 11023 12828 11176
rect 12894 11023 12904 11176
rect 13010 11023 13020 11176
rect 13086 11023 13096 11176
rect 13202 11023 13212 11176
rect 13278 11023 13288 11176
rect 13394 11023 13404 11176
rect 13470 11023 13480 11176
rect 13586 11023 13596 11176
rect 13662 11023 13672 11176
rect 13778 11023 13788 11176
rect 13854 11023 13864 11176
rect 13970 11023 13980 11176
rect 14046 11023 14056 11176
rect 14162 11023 14172 11176
rect 14238 11023 14248 11176
rect 14284 10963 14504 11210
rect 14646 11023 14656 11176
rect 14722 11023 14732 11176
rect 14838 11023 14848 11176
rect 14914 11023 14924 11176
rect 15030 11023 15040 11176
rect 15106 11023 15116 11176
rect 15222 11023 15232 11176
rect 15298 11023 15308 11176
rect 15414 11023 15424 11176
rect 15490 11023 15500 11176
rect 15606 11023 15616 11176
rect 15682 11023 15692 11176
rect 15798 11023 15808 11176
rect 15874 11023 15884 11176
rect 15990 11023 16000 11176
rect 16066 11023 16076 11176
rect 16112 10963 16332 11210
rect 16474 11023 16484 11176
rect 16550 11023 16560 11176
rect 16666 11023 16676 11176
rect 16742 11023 16752 11176
rect 16858 11023 16868 11176
rect 16934 11023 16944 11176
rect 17050 11023 17060 11176
rect 17126 11023 17136 11176
rect 17242 11023 17252 11176
rect 17318 11023 17328 11176
rect 17434 11023 17444 11176
rect 17510 11023 17520 11176
rect 17626 11023 17636 11176
rect 17702 11023 17712 11176
rect 17818 11023 17828 11176
rect 17894 11023 17904 11176
rect 17940 10963 18160 11210
rect 18302 11023 18312 11176
rect 18378 11023 18388 11176
rect 18494 11023 18504 11176
rect 18570 11023 18580 11176
rect 18686 11023 18696 11176
rect 18762 11023 18772 11176
rect 18878 11023 18888 11176
rect 18954 11023 18964 11176
rect 19070 11023 19080 11176
rect 19146 11023 19156 11176
rect 19262 11023 19272 11176
rect 19338 11023 19348 11176
rect 19454 11023 19464 11176
rect 19530 11023 19540 11176
rect 19646 11023 19656 11176
rect 19722 11023 19732 11176
rect 19768 10963 19988 11210
rect 20130 11023 20140 11176
rect 20206 11023 20216 11176
rect 20322 11023 20332 11176
rect 20398 11023 20408 11176
rect 20514 11023 20524 11176
rect 20590 11023 20600 11176
rect 20706 11023 20716 11176
rect 20782 11023 20792 11176
rect 20898 11023 20908 11176
rect 20974 11023 20984 11176
rect 21090 11023 21100 11176
rect 21166 11023 21176 11176
rect 21282 11023 21292 11176
rect 21358 11023 21368 11176
rect 21474 11023 21484 11176
rect 21550 11023 21560 11176
rect 21596 10963 21816 11210
rect 118 10810 128 10963
rect 194 10810 204 10963
rect 310 10810 320 10963
rect 386 10810 396 10963
rect 502 10810 512 10963
rect 578 10810 588 10963
rect 694 10810 704 10963
rect 770 10810 780 10963
rect 886 10810 896 10963
rect 962 10810 972 10963
rect 1078 10810 1088 10963
rect 1154 10810 1164 10963
rect 1270 10810 1280 10963
rect 1346 10810 1356 10963
rect 1462 10810 1472 10963
rect 1528 10810 1708 10963
rect 1946 10810 1956 10963
rect 2022 10810 2032 10963
rect 2138 10810 2148 10963
rect 2214 10810 2224 10963
rect 2330 10810 2340 10963
rect 2406 10810 2416 10963
rect 2522 10810 2532 10963
rect 2598 10810 2608 10963
rect 2714 10810 2724 10963
rect 2790 10810 2800 10963
rect 2906 10810 2916 10963
rect 2982 10810 2992 10963
rect 3098 10810 3108 10963
rect 3174 10810 3184 10963
rect 3290 10810 3300 10963
rect 3356 10810 3536 10963
rect 3774 10810 3784 10963
rect 3850 10810 3860 10963
rect 3966 10810 3976 10963
rect 4042 10810 4052 10963
rect 4158 10810 4168 10963
rect 4234 10810 4244 10963
rect 4350 10810 4360 10963
rect 4426 10810 4436 10963
rect 4542 10810 4552 10963
rect 4618 10810 4628 10963
rect 4734 10810 4744 10963
rect 4810 10810 4820 10963
rect 4926 10810 4936 10963
rect 5002 10810 5012 10963
rect 5118 10810 5128 10963
rect 5184 10810 5364 10963
rect 5602 10810 5612 10963
rect 5678 10810 5688 10963
rect 5794 10810 5804 10963
rect 5870 10810 5880 10963
rect 5986 10810 5996 10963
rect 6062 10810 6072 10963
rect 6178 10810 6188 10963
rect 6254 10810 6264 10963
rect 6370 10810 6380 10963
rect 6446 10810 6456 10963
rect 6562 10810 6572 10963
rect 6638 10810 6648 10963
rect 6754 10810 6764 10963
rect 6830 10810 6840 10963
rect 6946 10810 6956 10963
rect 7012 10810 7192 10963
rect 7430 10810 7440 10963
rect 7506 10810 7516 10963
rect 7622 10810 7632 10963
rect 7698 10810 7708 10963
rect 7814 10810 7824 10963
rect 7890 10810 7900 10963
rect 8006 10810 8016 10963
rect 8082 10810 8092 10963
rect 8198 10810 8208 10963
rect 8274 10810 8284 10963
rect 8390 10810 8400 10963
rect 8466 10810 8476 10963
rect 8582 10810 8592 10963
rect 8658 10810 8668 10963
rect 8774 10810 8784 10963
rect 8840 10810 9020 10963
rect 9258 10810 9268 10963
rect 9334 10810 9344 10963
rect 9450 10810 9460 10963
rect 9526 10810 9536 10963
rect 9642 10810 9652 10963
rect 9718 10810 9728 10963
rect 9834 10810 9844 10963
rect 9910 10810 9920 10963
rect 10026 10810 10036 10963
rect 10102 10810 10112 10963
rect 10218 10810 10228 10963
rect 10294 10810 10304 10963
rect 10410 10810 10420 10963
rect 10486 10810 10496 10963
rect 10602 10810 10612 10963
rect 10668 10810 10848 10963
rect 11086 10810 11096 10963
rect 11162 10810 11172 10963
rect 11278 10810 11288 10963
rect 11354 10810 11364 10963
rect 11470 10810 11480 10963
rect 11546 10810 11556 10963
rect 11662 10810 11672 10963
rect 11738 10810 11748 10963
rect 11854 10810 11864 10963
rect 11930 10810 11940 10963
rect 12046 10810 12056 10963
rect 12122 10810 12132 10963
rect 12238 10810 12248 10963
rect 12314 10810 12324 10963
rect 12430 10810 12440 10963
rect 12496 10810 12676 10963
rect 12914 10810 12924 10963
rect 12990 10810 13000 10963
rect 13106 10810 13116 10963
rect 13182 10810 13192 10963
rect 13298 10810 13308 10963
rect 13374 10810 13384 10963
rect 13490 10810 13500 10963
rect 13566 10810 13576 10963
rect 13682 10810 13692 10963
rect 13758 10810 13768 10963
rect 13874 10810 13884 10963
rect 13950 10810 13960 10963
rect 14066 10810 14076 10963
rect 14142 10810 14152 10963
rect 14258 10810 14268 10963
rect 14324 10810 14504 10963
rect 14742 10810 14752 10963
rect 14818 10810 14828 10963
rect 14934 10810 14944 10963
rect 15010 10810 15020 10963
rect 15126 10810 15136 10963
rect 15202 10810 15212 10963
rect 15318 10810 15328 10963
rect 15394 10810 15404 10963
rect 15510 10810 15520 10963
rect 15586 10810 15596 10963
rect 15702 10810 15712 10963
rect 15778 10810 15788 10963
rect 15894 10810 15904 10963
rect 15970 10810 15980 10963
rect 16086 10810 16096 10963
rect 16152 10810 16332 10963
rect 16570 10810 16580 10963
rect 16646 10810 16656 10963
rect 16762 10810 16772 10963
rect 16838 10810 16848 10963
rect 16954 10810 16964 10963
rect 17030 10810 17040 10963
rect 17146 10810 17156 10963
rect 17222 10810 17232 10963
rect 17338 10810 17348 10963
rect 17414 10810 17424 10963
rect 17530 10810 17540 10963
rect 17606 10810 17616 10963
rect 17722 10810 17732 10963
rect 17798 10810 17808 10963
rect 17914 10810 17924 10963
rect 17980 10810 18160 10963
rect 18398 10810 18408 10963
rect 18474 10810 18484 10963
rect 18590 10810 18600 10963
rect 18666 10810 18676 10963
rect 18782 10810 18792 10963
rect 18858 10810 18868 10963
rect 18974 10810 18984 10963
rect 19050 10810 19060 10963
rect 19166 10810 19176 10963
rect 19242 10810 19252 10963
rect 19358 10810 19368 10963
rect 19434 10810 19444 10963
rect 19550 10810 19560 10963
rect 19626 10810 19636 10963
rect 19742 10810 19752 10963
rect 19808 10810 19988 10963
rect 20226 10810 20236 10963
rect 20302 10810 20312 10963
rect 20418 10810 20428 10963
rect 20494 10810 20504 10963
rect 20610 10810 20620 10963
rect 20686 10810 20696 10963
rect 20802 10810 20812 10963
rect 20878 10810 20888 10963
rect 20994 10810 21004 10963
rect 21070 10810 21080 10963
rect 21186 10810 21196 10963
rect 21262 10810 21272 10963
rect 21378 10810 21388 10963
rect 21454 10810 21464 10963
rect 21570 10810 21580 10963
rect 21636 10810 21816 10963
rect 0 10713 1490 10772
rect 1828 10713 3318 10772
rect 3656 10713 5146 10772
rect 5484 10713 6974 10772
rect 7312 10713 8802 10772
rect 9140 10713 10630 10772
rect 10968 10713 12458 10772
rect 12796 10713 14286 10772
rect 14624 10713 16114 10772
rect 16452 10713 17942 10772
rect 18280 10713 19770 10772
rect 20108 10713 21598 10772
rect 0 10534 1490 10593
rect 1828 10534 3318 10593
rect 3656 10534 5146 10593
rect 5484 10534 6974 10593
rect 7312 10534 8802 10593
rect 9140 10534 10630 10593
rect 10968 10534 12458 10593
rect 12796 10534 14286 10593
rect 14624 10534 16114 10593
rect 16452 10534 17942 10593
rect 18280 10534 19770 10593
rect 20108 10534 21598 10593
rect 22 10309 32 10462
rect 98 10309 108 10462
rect 214 10309 224 10462
rect 290 10309 300 10462
rect 406 10309 416 10462
rect 482 10309 492 10462
rect 598 10309 608 10462
rect 674 10309 684 10462
rect 790 10309 800 10462
rect 866 10309 876 10462
rect 982 10309 992 10462
rect 1058 10309 1068 10462
rect 1174 10309 1184 10462
rect 1250 10309 1260 10462
rect 1366 10309 1376 10462
rect 1442 10309 1452 10462
rect 1488 10249 1708 10496
rect 1850 10309 1860 10462
rect 1926 10309 1936 10462
rect 2042 10309 2052 10462
rect 2118 10309 2128 10462
rect 2234 10309 2244 10462
rect 2310 10309 2320 10462
rect 2426 10309 2436 10462
rect 2502 10309 2512 10462
rect 2618 10309 2628 10462
rect 2694 10309 2704 10462
rect 2810 10309 2820 10462
rect 2886 10309 2896 10462
rect 3002 10309 3012 10462
rect 3078 10309 3088 10462
rect 3194 10309 3204 10462
rect 3270 10309 3280 10462
rect 3316 10249 3536 10496
rect 3678 10309 3688 10462
rect 3754 10309 3764 10462
rect 3870 10309 3880 10462
rect 3946 10309 3956 10462
rect 4062 10309 4072 10462
rect 4138 10309 4148 10462
rect 4254 10309 4264 10462
rect 4330 10309 4340 10462
rect 4446 10309 4456 10462
rect 4522 10309 4532 10462
rect 4638 10309 4648 10462
rect 4714 10309 4724 10462
rect 4830 10309 4840 10462
rect 4906 10309 4916 10462
rect 5022 10309 5032 10462
rect 5098 10309 5108 10462
rect 5144 10249 5364 10496
rect 5506 10309 5516 10462
rect 5582 10309 5592 10462
rect 5698 10309 5708 10462
rect 5774 10309 5784 10462
rect 5890 10309 5900 10462
rect 5966 10309 5976 10462
rect 6082 10309 6092 10462
rect 6158 10309 6168 10462
rect 6274 10309 6284 10462
rect 6350 10309 6360 10462
rect 6466 10309 6476 10462
rect 6542 10309 6552 10462
rect 6658 10309 6668 10462
rect 6734 10309 6744 10462
rect 6850 10309 6860 10462
rect 6926 10309 6936 10462
rect 6972 10249 7192 10496
rect 7334 10309 7344 10462
rect 7410 10309 7420 10462
rect 7526 10309 7536 10462
rect 7602 10309 7612 10462
rect 7718 10309 7728 10462
rect 7794 10309 7804 10462
rect 7910 10309 7920 10462
rect 7986 10309 7996 10462
rect 8102 10309 8112 10462
rect 8178 10309 8188 10462
rect 8294 10309 8304 10462
rect 8370 10309 8380 10462
rect 8486 10309 8496 10462
rect 8562 10309 8572 10462
rect 8678 10309 8688 10462
rect 8754 10309 8764 10462
rect 8800 10249 9020 10496
rect 9162 10309 9172 10462
rect 9238 10309 9248 10462
rect 9354 10309 9364 10462
rect 9430 10309 9440 10462
rect 9546 10309 9556 10462
rect 9622 10309 9632 10462
rect 9738 10309 9748 10462
rect 9814 10309 9824 10462
rect 9930 10309 9940 10462
rect 10006 10309 10016 10462
rect 10122 10309 10132 10462
rect 10198 10309 10208 10462
rect 10314 10309 10324 10462
rect 10390 10309 10400 10462
rect 10506 10309 10516 10462
rect 10582 10309 10592 10462
rect 10628 10249 10848 10496
rect 10990 10309 11000 10462
rect 11066 10309 11076 10462
rect 11182 10309 11192 10462
rect 11258 10309 11268 10462
rect 11374 10309 11384 10462
rect 11450 10309 11460 10462
rect 11566 10309 11576 10462
rect 11642 10309 11652 10462
rect 11758 10309 11768 10462
rect 11834 10309 11844 10462
rect 11950 10309 11960 10462
rect 12026 10309 12036 10462
rect 12142 10309 12152 10462
rect 12218 10309 12228 10462
rect 12334 10309 12344 10462
rect 12410 10309 12420 10462
rect 12456 10249 12676 10496
rect 12818 10309 12828 10462
rect 12894 10309 12904 10462
rect 13010 10309 13020 10462
rect 13086 10309 13096 10462
rect 13202 10309 13212 10462
rect 13278 10309 13288 10462
rect 13394 10309 13404 10462
rect 13470 10309 13480 10462
rect 13586 10309 13596 10462
rect 13662 10309 13672 10462
rect 13778 10309 13788 10462
rect 13854 10309 13864 10462
rect 13970 10309 13980 10462
rect 14046 10309 14056 10462
rect 14162 10309 14172 10462
rect 14238 10309 14248 10462
rect 14284 10249 14504 10496
rect 14646 10309 14656 10462
rect 14722 10309 14732 10462
rect 14838 10309 14848 10462
rect 14914 10309 14924 10462
rect 15030 10309 15040 10462
rect 15106 10309 15116 10462
rect 15222 10309 15232 10462
rect 15298 10309 15308 10462
rect 15414 10309 15424 10462
rect 15490 10309 15500 10462
rect 15606 10309 15616 10462
rect 15682 10309 15692 10462
rect 15798 10309 15808 10462
rect 15874 10309 15884 10462
rect 15990 10309 16000 10462
rect 16066 10309 16076 10462
rect 16112 10249 16332 10496
rect 16474 10309 16484 10462
rect 16550 10309 16560 10462
rect 16666 10309 16676 10462
rect 16742 10309 16752 10462
rect 16858 10309 16868 10462
rect 16934 10309 16944 10462
rect 17050 10309 17060 10462
rect 17126 10309 17136 10462
rect 17242 10309 17252 10462
rect 17318 10309 17328 10462
rect 17434 10309 17444 10462
rect 17510 10309 17520 10462
rect 17626 10309 17636 10462
rect 17702 10309 17712 10462
rect 17818 10309 17828 10462
rect 17894 10309 17904 10462
rect 17940 10249 18160 10496
rect 18302 10309 18312 10462
rect 18378 10309 18388 10462
rect 18494 10309 18504 10462
rect 18570 10309 18580 10462
rect 18686 10309 18696 10462
rect 18762 10309 18772 10462
rect 18878 10309 18888 10462
rect 18954 10309 18964 10462
rect 19070 10309 19080 10462
rect 19146 10309 19156 10462
rect 19262 10309 19272 10462
rect 19338 10309 19348 10462
rect 19454 10309 19464 10462
rect 19530 10309 19540 10462
rect 19646 10309 19656 10462
rect 19722 10309 19732 10462
rect 19768 10249 19988 10496
rect 20130 10309 20140 10462
rect 20206 10309 20216 10462
rect 20322 10309 20332 10462
rect 20398 10309 20408 10462
rect 20514 10309 20524 10462
rect 20590 10309 20600 10462
rect 20706 10309 20716 10462
rect 20782 10309 20792 10462
rect 20898 10309 20908 10462
rect 20974 10309 20984 10462
rect 21090 10309 21100 10462
rect 21166 10309 21176 10462
rect 21282 10309 21292 10462
rect 21358 10309 21368 10462
rect 21474 10309 21484 10462
rect 21550 10309 21560 10462
rect 21596 10249 21816 10496
rect 118 10096 128 10249
rect 194 10096 204 10249
rect 310 10096 320 10249
rect 386 10096 396 10249
rect 502 10096 512 10249
rect 578 10096 588 10249
rect 694 10096 704 10249
rect 770 10096 780 10249
rect 886 10096 896 10249
rect 962 10096 972 10249
rect 1078 10096 1088 10249
rect 1154 10096 1164 10249
rect 1270 10096 1280 10249
rect 1346 10096 1356 10249
rect 1462 10096 1472 10249
rect 1528 10096 1708 10249
rect 1946 10096 1956 10249
rect 2022 10096 2032 10249
rect 2138 10096 2148 10249
rect 2214 10096 2224 10249
rect 2330 10096 2340 10249
rect 2406 10096 2416 10249
rect 2522 10096 2532 10249
rect 2598 10096 2608 10249
rect 2714 10096 2724 10249
rect 2790 10096 2800 10249
rect 2906 10096 2916 10249
rect 2982 10096 2992 10249
rect 3098 10096 3108 10249
rect 3174 10096 3184 10249
rect 3290 10096 3300 10249
rect 3356 10096 3536 10249
rect 3774 10096 3784 10249
rect 3850 10096 3860 10249
rect 3966 10096 3976 10249
rect 4042 10096 4052 10249
rect 4158 10096 4168 10249
rect 4234 10096 4244 10249
rect 4350 10096 4360 10249
rect 4426 10096 4436 10249
rect 4542 10096 4552 10249
rect 4618 10096 4628 10249
rect 4734 10096 4744 10249
rect 4810 10096 4820 10249
rect 4926 10096 4936 10249
rect 5002 10096 5012 10249
rect 5118 10096 5128 10249
rect 5184 10096 5364 10249
rect 5602 10096 5612 10249
rect 5678 10096 5688 10249
rect 5794 10096 5804 10249
rect 5870 10096 5880 10249
rect 5986 10096 5996 10249
rect 6062 10096 6072 10249
rect 6178 10096 6188 10249
rect 6254 10096 6264 10249
rect 6370 10096 6380 10249
rect 6446 10096 6456 10249
rect 6562 10096 6572 10249
rect 6638 10096 6648 10249
rect 6754 10096 6764 10249
rect 6830 10096 6840 10249
rect 6946 10096 6956 10249
rect 7012 10096 7192 10249
rect 7430 10096 7440 10249
rect 7506 10096 7516 10249
rect 7622 10096 7632 10249
rect 7698 10096 7708 10249
rect 7814 10096 7824 10249
rect 7890 10096 7900 10249
rect 8006 10096 8016 10249
rect 8082 10096 8092 10249
rect 8198 10096 8208 10249
rect 8274 10096 8284 10249
rect 8390 10096 8400 10249
rect 8466 10096 8476 10249
rect 8582 10096 8592 10249
rect 8658 10096 8668 10249
rect 8774 10096 8784 10249
rect 8840 10096 9020 10249
rect 9258 10096 9268 10249
rect 9334 10096 9344 10249
rect 9450 10096 9460 10249
rect 9526 10096 9536 10249
rect 9642 10096 9652 10249
rect 9718 10096 9728 10249
rect 9834 10096 9844 10249
rect 9910 10096 9920 10249
rect 10026 10096 10036 10249
rect 10102 10096 10112 10249
rect 10218 10096 10228 10249
rect 10294 10096 10304 10249
rect 10410 10096 10420 10249
rect 10486 10096 10496 10249
rect 10602 10096 10612 10249
rect 10668 10096 10848 10249
rect 11086 10096 11096 10249
rect 11162 10096 11172 10249
rect 11278 10096 11288 10249
rect 11354 10096 11364 10249
rect 11470 10096 11480 10249
rect 11546 10096 11556 10249
rect 11662 10096 11672 10249
rect 11738 10096 11748 10249
rect 11854 10096 11864 10249
rect 11930 10096 11940 10249
rect 12046 10096 12056 10249
rect 12122 10096 12132 10249
rect 12238 10096 12248 10249
rect 12314 10096 12324 10249
rect 12430 10096 12440 10249
rect 12496 10096 12676 10249
rect 12914 10096 12924 10249
rect 12990 10096 13000 10249
rect 13106 10096 13116 10249
rect 13182 10096 13192 10249
rect 13298 10096 13308 10249
rect 13374 10096 13384 10249
rect 13490 10096 13500 10249
rect 13566 10096 13576 10249
rect 13682 10096 13692 10249
rect 13758 10096 13768 10249
rect 13874 10096 13884 10249
rect 13950 10096 13960 10249
rect 14066 10096 14076 10249
rect 14142 10096 14152 10249
rect 14258 10096 14268 10249
rect 14324 10096 14504 10249
rect 14742 10096 14752 10249
rect 14818 10096 14828 10249
rect 14934 10096 14944 10249
rect 15010 10096 15020 10249
rect 15126 10096 15136 10249
rect 15202 10096 15212 10249
rect 15318 10096 15328 10249
rect 15394 10096 15404 10249
rect 15510 10096 15520 10249
rect 15586 10096 15596 10249
rect 15702 10096 15712 10249
rect 15778 10096 15788 10249
rect 15894 10096 15904 10249
rect 15970 10096 15980 10249
rect 16086 10096 16096 10249
rect 16152 10096 16332 10249
rect 16570 10096 16580 10249
rect 16646 10096 16656 10249
rect 16762 10096 16772 10249
rect 16838 10096 16848 10249
rect 16954 10096 16964 10249
rect 17030 10096 17040 10249
rect 17146 10096 17156 10249
rect 17222 10096 17232 10249
rect 17338 10096 17348 10249
rect 17414 10096 17424 10249
rect 17530 10096 17540 10249
rect 17606 10096 17616 10249
rect 17722 10096 17732 10249
rect 17798 10096 17808 10249
rect 17914 10096 17924 10249
rect 17980 10096 18160 10249
rect 18398 10096 18408 10249
rect 18474 10096 18484 10249
rect 18590 10096 18600 10249
rect 18666 10096 18676 10249
rect 18782 10096 18792 10249
rect 18858 10096 18868 10249
rect 18974 10096 18984 10249
rect 19050 10096 19060 10249
rect 19166 10096 19176 10249
rect 19242 10096 19252 10249
rect 19358 10096 19368 10249
rect 19434 10096 19444 10249
rect 19550 10096 19560 10249
rect 19626 10096 19636 10249
rect 19742 10096 19752 10249
rect 19808 10096 19988 10249
rect 20226 10096 20236 10249
rect 20302 10096 20312 10249
rect 20418 10096 20428 10249
rect 20494 10096 20504 10249
rect 20610 10096 20620 10249
rect 20686 10096 20696 10249
rect 20802 10096 20812 10249
rect 20878 10096 20888 10249
rect 20994 10096 21004 10249
rect 21070 10096 21080 10249
rect 21186 10096 21196 10249
rect 21262 10096 21272 10249
rect 21378 10096 21388 10249
rect 21454 10096 21464 10249
rect 21570 10096 21580 10249
rect 21636 10096 21816 10249
rect 0 9999 1490 10058
rect 1828 9999 3318 10058
rect 3656 9999 5146 10058
rect 5484 9999 6974 10058
rect 7312 9999 8802 10058
rect 9140 9999 10630 10058
rect 10968 9999 12458 10058
rect 12796 9999 14286 10058
rect 14624 9999 16114 10058
rect 16452 9999 17942 10058
rect 18280 9999 19770 10058
rect 20108 9999 21598 10058
rect 0 9820 1490 9879
rect 1828 9820 3318 9879
rect 3656 9820 5146 9879
rect 5484 9820 6974 9879
rect 7312 9820 8802 9879
rect 9140 9820 10630 9879
rect 10968 9820 12458 9879
rect 12796 9820 14286 9879
rect 14624 9820 16114 9879
rect 16452 9820 17942 9879
rect 18280 9820 19770 9879
rect 20108 9820 21598 9879
rect 22 9595 32 9748
rect 98 9595 108 9748
rect 214 9595 224 9748
rect 290 9595 300 9748
rect 406 9595 416 9748
rect 482 9595 492 9748
rect 598 9595 608 9748
rect 674 9595 684 9748
rect 790 9595 800 9748
rect 866 9595 876 9748
rect 982 9595 992 9748
rect 1058 9595 1068 9748
rect 1174 9595 1184 9748
rect 1250 9595 1260 9748
rect 1366 9595 1376 9748
rect 1442 9595 1452 9748
rect 1488 9535 1708 9782
rect 1850 9595 1860 9748
rect 1926 9595 1936 9748
rect 2042 9595 2052 9748
rect 2118 9595 2128 9748
rect 2234 9595 2244 9748
rect 2310 9595 2320 9748
rect 2426 9595 2436 9748
rect 2502 9595 2512 9748
rect 2618 9595 2628 9748
rect 2694 9595 2704 9748
rect 2810 9595 2820 9748
rect 2886 9595 2896 9748
rect 3002 9595 3012 9748
rect 3078 9595 3088 9748
rect 3194 9595 3204 9748
rect 3270 9595 3280 9748
rect 3316 9535 3536 9782
rect 3678 9595 3688 9748
rect 3754 9595 3764 9748
rect 3870 9595 3880 9748
rect 3946 9595 3956 9748
rect 4062 9595 4072 9748
rect 4138 9595 4148 9748
rect 4254 9595 4264 9748
rect 4330 9595 4340 9748
rect 4446 9595 4456 9748
rect 4522 9595 4532 9748
rect 4638 9595 4648 9748
rect 4714 9595 4724 9748
rect 4830 9595 4840 9748
rect 4906 9595 4916 9748
rect 5022 9595 5032 9748
rect 5098 9595 5108 9748
rect 5144 9535 5364 9782
rect 5506 9595 5516 9748
rect 5582 9595 5592 9748
rect 5698 9595 5708 9748
rect 5774 9595 5784 9748
rect 5890 9595 5900 9748
rect 5966 9595 5976 9748
rect 6082 9595 6092 9748
rect 6158 9595 6168 9748
rect 6274 9595 6284 9748
rect 6350 9595 6360 9748
rect 6466 9595 6476 9748
rect 6542 9595 6552 9748
rect 6658 9595 6668 9748
rect 6734 9595 6744 9748
rect 6850 9595 6860 9748
rect 6926 9595 6936 9748
rect 6972 9535 7192 9782
rect 7334 9595 7344 9748
rect 7410 9595 7420 9748
rect 7526 9595 7536 9748
rect 7602 9595 7612 9748
rect 7718 9595 7728 9748
rect 7794 9595 7804 9748
rect 7910 9595 7920 9748
rect 7986 9595 7996 9748
rect 8102 9595 8112 9748
rect 8178 9595 8188 9748
rect 8294 9595 8304 9748
rect 8370 9595 8380 9748
rect 8486 9595 8496 9748
rect 8562 9595 8572 9748
rect 8678 9595 8688 9748
rect 8754 9595 8764 9748
rect 8800 9535 9020 9782
rect 9162 9595 9172 9748
rect 9238 9595 9248 9748
rect 9354 9595 9364 9748
rect 9430 9595 9440 9748
rect 9546 9595 9556 9748
rect 9622 9595 9632 9748
rect 9738 9595 9748 9748
rect 9814 9595 9824 9748
rect 9930 9595 9940 9748
rect 10006 9595 10016 9748
rect 10122 9595 10132 9748
rect 10198 9595 10208 9748
rect 10314 9595 10324 9748
rect 10390 9595 10400 9748
rect 10506 9595 10516 9748
rect 10582 9595 10592 9748
rect 10628 9535 10848 9782
rect 10990 9595 11000 9748
rect 11066 9595 11076 9748
rect 11182 9595 11192 9748
rect 11258 9595 11268 9748
rect 11374 9595 11384 9748
rect 11450 9595 11460 9748
rect 11566 9595 11576 9748
rect 11642 9595 11652 9748
rect 11758 9595 11768 9748
rect 11834 9595 11844 9748
rect 11950 9595 11960 9748
rect 12026 9595 12036 9748
rect 12142 9595 12152 9748
rect 12218 9595 12228 9748
rect 12334 9595 12344 9748
rect 12410 9595 12420 9748
rect 12456 9535 12676 9782
rect 12818 9595 12828 9748
rect 12894 9595 12904 9748
rect 13010 9595 13020 9748
rect 13086 9595 13096 9748
rect 13202 9595 13212 9748
rect 13278 9595 13288 9748
rect 13394 9595 13404 9748
rect 13470 9595 13480 9748
rect 13586 9595 13596 9748
rect 13662 9595 13672 9748
rect 13778 9595 13788 9748
rect 13854 9595 13864 9748
rect 13970 9595 13980 9748
rect 14046 9595 14056 9748
rect 14162 9595 14172 9748
rect 14238 9595 14248 9748
rect 14284 9535 14504 9782
rect 14646 9595 14656 9748
rect 14722 9595 14732 9748
rect 14838 9595 14848 9748
rect 14914 9595 14924 9748
rect 15030 9595 15040 9748
rect 15106 9595 15116 9748
rect 15222 9595 15232 9748
rect 15298 9595 15308 9748
rect 15414 9595 15424 9748
rect 15490 9595 15500 9748
rect 15606 9595 15616 9748
rect 15682 9595 15692 9748
rect 15798 9595 15808 9748
rect 15874 9595 15884 9748
rect 15990 9595 16000 9748
rect 16066 9595 16076 9748
rect 16112 9535 16332 9782
rect 16474 9595 16484 9748
rect 16550 9595 16560 9748
rect 16666 9595 16676 9748
rect 16742 9595 16752 9748
rect 16858 9595 16868 9748
rect 16934 9595 16944 9748
rect 17050 9595 17060 9748
rect 17126 9595 17136 9748
rect 17242 9595 17252 9748
rect 17318 9595 17328 9748
rect 17434 9595 17444 9748
rect 17510 9595 17520 9748
rect 17626 9595 17636 9748
rect 17702 9595 17712 9748
rect 17818 9595 17828 9748
rect 17894 9595 17904 9748
rect 17940 9535 18160 9782
rect 18302 9595 18312 9748
rect 18378 9595 18388 9748
rect 18494 9595 18504 9748
rect 18570 9595 18580 9748
rect 18686 9595 18696 9748
rect 18762 9595 18772 9748
rect 18878 9595 18888 9748
rect 18954 9595 18964 9748
rect 19070 9595 19080 9748
rect 19146 9595 19156 9748
rect 19262 9595 19272 9748
rect 19338 9595 19348 9748
rect 19454 9595 19464 9748
rect 19530 9595 19540 9748
rect 19646 9595 19656 9748
rect 19722 9595 19732 9748
rect 19768 9535 19988 9782
rect 20130 9595 20140 9748
rect 20206 9595 20216 9748
rect 20322 9595 20332 9748
rect 20398 9595 20408 9748
rect 20514 9595 20524 9748
rect 20590 9595 20600 9748
rect 20706 9595 20716 9748
rect 20782 9595 20792 9748
rect 20898 9595 20908 9748
rect 20974 9595 20984 9748
rect 21090 9595 21100 9748
rect 21166 9595 21176 9748
rect 21282 9595 21292 9748
rect 21358 9595 21368 9748
rect 21474 9595 21484 9748
rect 21550 9595 21560 9748
rect 21596 9535 21816 9782
rect 118 9382 128 9535
rect 194 9382 204 9535
rect 310 9382 320 9535
rect 386 9382 396 9535
rect 502 9382 512 9535
rect 578 9382 588 9535
rect 694 9382 704 9535
rect 770 9382 780 9535
rect 886 9382 896 9535
rect 962 9382 972 9535
rect 1078 9382 1088 9535
rect 1154 9382 1164 9535
rect 1270 9382 1280 9535
rect 1346 9382 1356 9535
rect 1462 9382 1472 9535
rect 1528 9382 1708 9535
rect 1946 9382 1956 9535
rect 2022 9382 2032 9535
rect 2138 9382 2148 9535
rect 2214 9382 2224 9535
rect 2330 9382 2340 9535
rect 2406 9382 2416 9535
rect 2522 9382 2532 9535
rect 2598 9382 2608 9535
rect 2714 9382 2724 9535
rect 2790 9382 2800 9535
rect 2906 9382 2916 9535
rect 2982 9382 2992 9535
rect 3098 9382 3108 9535
rect 3174 9382 3184 9535
rect 3290 9382 3300 9535
rect 3356 9382 3536 9535
rect 3774 9382 3784 9535
rect 3850 9382 3860 9535
rect 3966 9382 3976 9535
rect 4042 9382 4052 9535
rect 4158 9382 4168 9535
rect 4234 9382 4244 9535
rect 4350 9382 4360 9535
rect 4426 9382 4436 9535
rect 4542 9382 4552 9535
rect 4618 9382 4628 9535
rect 4734 9382 4744 9535
rect 4810 9382 4820 9535
rect 4926 9382 4936 9535
rect 5002 9382 5012 9535
rect 5118 9382 5128 9535
rect 5184 9382 5364 9535
rect 5602 9382 5612 9535
rect 5678 9382 5688 9535
rect 5794 9382 5804 9535
rect 5870 9382 5880 9535
rect 5986 9382 5996 9535
rect 6062 9382 6072 9535
rect 6178 9382 6188 9535
rect 6254 9382 6264 9535
rect 6370 9382 6380 9535
rect 6446 9382 6456 9535
rect 6562 9382 6572 9535
rect 6638 9382 6648 9535
rect 6754 9382 6764 9535
rect 6830 9382 6840 9535
rect 6946 9382 6956 9535
rect 7012 9382 7192 9535
rect 7430 9382 7440 9535
rect 7506 9382 7516 9535
rect 7622 9382 7632 9535
rect 7698 9382 7708 9535
rect 7814 9382 7824 9535
rect 7890 9382 7900 9535
rect 8006 9382 8016 9535
rect 8082 9382 8092 9535
rect 8198 9382 8208 9535
rect 8274 9382 8284 9535
rect 8390 9382 8400 9535
rect 8466 9382 8476 9535
rect 8582 9382 8592 9535
rect 8658 9382 8668 9535
rect 8774 9382 8784 9535
rect 8840 9382 9020 9535
rect 9258 9382 9268 9535
rect 9334 9382 9344 9535
rect 9450 9382 9460 9535
rect 9526 9382 9536 9535
rect 9642 9382 9652 9535
rect 9718 9382 9728 9535
rect 9834 9382 9844 9535
rect 9910 9382 9920 9535
rect 10026 9382 10036 9535
rect 10102 9382 10112 9535
rect 10218 9382 10228 9535
rect 10294 9382 10304 9535
rect 10410 9382 10420 9535
rect 10486 9382 10496 9535
rect 10602 9382 10612 9535
rect 10668 9382 10848 9535
rect 11086 9382 11096 9535
rect 11162 9382 11172 9535
rect 11278 9382 11288 9535
rect 11354 9382 11364 9535
rect 11470 9382 11480 9535
rect 11546 9382 11556 9535
rect 11662 9382 11672 9535
rect 11738 9382 11748 9535
rect 11854 9382 11864 9535
rect 11930 9382 11940 9535
rect 12046 9382 12056 9535
rect 12122 9382 12132 9535
rect 12238 9382 12248 9535
rect 12314 9382 12324 9535
rect 12430 9382 12440 9535
rect 12496 9382 12676 9535
rect 12914 9382 12924 9535
rect 12990 9382 13000 9535
rect 13106 9382 13116 9535
rect 13182 9382 13192 9535
rect 13298 9382 13308 9535
rect 13374 9382 13384 9535
rect 13490 9382 13500 9535
rect 13566 9382 13576 9535
rect 13682 9382 13692 9535
rect 13758 9382 13768 9535
rect 13874 9382 13884 9535
rect 13950 9382 13960 9535
rect 14066 9382 14076 9535
rect 14142 9382 14152 9535
rect 14258 9382 14268 9535
rect 14324 9382 14504 9535
rect 14742 9382 14752 9535
rect 14818 9382 14828 9535
rect 14934 9382 14944 9535
rect 15010 9382 15020 9535
rect 15126 9382 15136 9535
rect 15202 9382 15212 9535
rect 15318 9382 15328 9535
rect 15394 9382 15404 9535
rect 15510 9382 15520 9535
rect 15586 9382 15596 9535
rect 15702 9382 15712 9535
rect 15778 9382 15788 9535
rect 15894 9382 15904 9535
rect 15970 9382 15980 9535
rect 16086 9382 16096 9535
rect 16152 9382 16332 9535
rect 16570 9382 16580 9535
rect 16646 9382 16656 9535
rect 16762 9382 16772 9535
rect 16838 9382 16848 9535
rect 16954 9382 16964 9535
rect 17030 9382 17040 9535
rect 17146 9382 17156 9535
rect 17222 9382 17232 9535
rect 17338 9382 17348 9535
rect 17414 9382 17424 9535
rect 17530 9382 17540 9535
rect 17606 9382 17616 9535
rect 17722 9382 17732 9535
rect 17798 9382 17808 9535
rect 17914 9382 17924 9535
rect 17980 9382 18160 9535
rect 18398 9382 18408 9535
rect 18474 9382 18484 9535
rect 18590 9382 18600 9535
rect 18666 9382 18676 9535
rect 18782 9382 18792 9535
rect 18858 9382 18868 9535
rect 18974 9382 18984 9535
rect 19050 9382 19060 9535
rect 19166 9382 19176 9535
rect 19242 9382 19252 9535
rect 19358 9382 19368 9535
rect 19434 9382 19444 9535
rect 19550 9382 19560 9535
rect 19626 9382 19636 9535
rect 19742 9382 19752 9535
rect 19808 9382 19988 9535
rect 20226 9382 20236 9535
rect 20302 9382 20312 9535
rect 20418 9382 20428 9535
rect 20494 9382 20504 9535
rect 20610 9382 20620 9535
rect 20686 9382 20696 9535
rect 20802 9382 20812 9535
rect 20878 9382 20888 9535
rect 20994 9382 21004 9535
rect 21070 9382 21080 9535
rect 21186 9382 21196 9535
rect 21262 9382 21272 9535
rect 21378 9382 21388 9535
rect 21454 9382 21464 9535
rect 21570 9382 21580 9535
rect 21636 9382 21816 9535
rect 0 9285 1490 9344
rect 1828 9285 3318 9344
rect 3656 9285 5146 9344
rect 5484 9285 6974 9344
rect 7312 9285 8802 9344
rect 9140 9285 10630 9344
rect 10968 9285 12458 9344
rect 12796 9285 14286 9344
rect 14624 9285 16114 9344
rect 16452 9285 17942 9344
rect 18280 9285 19770 9344
rect 20108 9285 21598 9344
rect 0 9106 1490 9165
rect 1828 9106 3318 9165
rect 3656 9106 5146 9165
rect 5484 9106 6974 9165
rect 7312 9106 8802 9165
rect 9140 9106 10630 9165
rect 10968 9106 12458 9165
rect 12796 9106 14286 9165
rect 14624 9106 16114 9165
rect 16452 9106 17942 9165
rect 18280 9106 19770 9165
rect 20108 9106 21598 9165
rect 22 8881 32 9034
rect 98 8881 108 9034
rect 214 8881 224 9034
rect 290 8881 300 9034
rect 406 8881 416 9034
rect 482 8881 492 9034
rect 598 8881 608 9034
rect 674 8881 684 9034
rect 790 8881 800 9034
rect 866 8881 876 9034
rect 982 8881 992 9034
rect 1058 8881 1068 9034
rect 1174 8881 1184 9034
rect 1250 8881 1260 9034
rect 1366 8881 1376 9034
rect 1442 8881 1452 9034
rect 1488 8821 1708 9068
rect 1850 8881 1860 9034
rect 1926 8881 1936 9034
rect 2042 8881 2052 9034
rect 2118 8881 2128 9034
rect 2234 8881 2244 9034
rect 2310 8881 2320 9034
rect 2426 8881 2436 9034
rect 2502 8881 2512 9034
rect 2618 8881 2628 9034
rect 2694 8881 2704 9034
rect 2810 8881 2820 9034
rect 2886 8881 2896 9034
rect 3002 8881 3012 9034
rect 3078 8881 3088 9034
rect 3194 8881 3204 9034
rect 3270 8881 3280 9034
rect 3316 8821 3536 9068
rect 3678 8881 3688 9034
rect 3754 8881 3764 9034
rect 3870 8881 3880 9034
rect 3946 8881 3956 9034
rect 4062 8881 4072 9034
rect 4138 8881 4148 9034
rect 4254 8881 4264 9034
rect 4330 8881 4340 9034
rect 4446 8881 4456 9034
rect 4522 8881 4532 9034
rect 4638 8881 4648 9034
rect 4714 8881 4724 9034
rect 4830 8881 4840 9034
rect 4906 8881 4916 9034
rect 5022 8881 5032 9034
rect 5098 8881 5108 9034
rect 5144 8821 5364 9068
rect 5506 8881 5516 9034
rect 5582 8881 5592 9034
rect 5698 8881 5708 9034
rect 5774 8881 5784 9034
rect 5890 8881 5900 9034
rect 5966 8881 5976 9034
rect 6082 8881 6092 9034
rect 6158 8881 6168 9034
rect 6274 8881 6284 9034
rect 6350 8881 6360 9034
rect 6466 8881 6476 9034
rect 6542 8881 6552 9034
rect 6658 8881 6668 9034
rect 6734 8881 6744 9034
rect 6850 8881 6860 9034
rect 6926 8881 6936 9034
rect 6972 8821 7192 9068
rect 7334 8881 7344 9034
rect 7410 8881 7420 9034
rect 7526 8881 7536 9034
rect 7602 8881 7612 9034
rect 7718 8881 7728 9034
rect 7794 8881 7804 9034
rect 7910 8881 7920 9034
rect 7986 8881 7996 9034
rect 8102 8881 8112 9034
rect 8178 8881 8188 9034
rect 8294 8881 8304 9034
rect 8370 8881 8380 9034
rect 8486 8881 8496 9034
rect 8562 8881 8572 9034
rect 8678 8881 8688 9034
rect 8754 8881 8764 9034
rect 8800 8821 9020 9068
rect 9162 8881 9172 9034
rect 9238 8881 9248 9034
rect 9354 8881 9364 9034
rect 9430 8881 9440 9034
rect 9546 8881 9556 9034
rect 9622 8881 9632 9034
rect 9738 8881 9748 9034
rect 9814 8881 9824 9034
rect 9930 8881 9940 9034
rect 10006 8881 10016 9034
rect 10122 8881 10132 9034
rect 10198 8881 10208 9034
rect 10314 8881 10324 9034
rect 10390 8881 10400 9034
rect 10506 8881 10516 9034
rect 10582 8881 10592 9034
rect 10628 8821 10848 9068
rect 10990 8881 11000 9034
rect 11066 8881 11076 9034
rect 11182 8881 11192 9034
rect 11258 8881 11268 9034
rect 11374 8881 11384 9034
rect 11450 8881 11460 9034
rect 11566 8881 11576 9034
rect 11642 8881 11652 9034
rect 11758 8881 11768 9034
rect 11834 8881 11844 9034
rect 11950 8881 11960 9034
rect 12026 8881 12036 9034
rect 12142 8881 12152 9034
rect 12218 8881 12228 9034
rect 12334 8881 12344 9034
rect 12410 8881 12420 9034
rect 12456 8821 12676 9068
rect 12818 8881 12828 9034
rect 12894 8881 12904 9034
rect 13010 8881 13020 9034
rect 13086 8881 13096 9034
rect 13202 8881 13212 9034
rect 13278 8881 13288 9034
rect 13394 8881 13404 9034
rect 13470 8881 13480 9034
rect 13586 8881 13596 9034
rect 13662 8881 13672 9034
rect 13778 8881 13788 9034
rect 13854 8881 13864 9034
rect 13970 8881 13980 9034
rect 14046 8881 14056 9034
rect 14162 8881 14172 9034
rect 14238 8881 14248 9034
rect 14284 8821 14504 9068
rect 14646 8881 14656 9034
rect 14722 8881 14732 9034
rect 14838 8881 14848 9034
rect 14914 8881 14924 9034
rect 15030 8881 15040 9034
rect 15106 8881 15116 9034
rect 15222 8881 15232 9034
rect 15298 8881 15308 9034
rect 15414 8881 15424 9034
rect 15490 8881 15500 9034
rect 15606 8881 15616 9034
rect 15682 8881 15692 9034
rect 15798 8881 15808 9034
rect 15874 8881 15884 9034
rect 15990 8881 16000 9034
rect 16066 8881 16076 9034
rect 16112 8821 16332 9068
rect 16474 8881 16484 9034
rect 16550 8881 16560 9034
rect 16666 8881 16676 9034
rect 16742 8881 16752 9034
rect 16858 8881 16868 9034
rect 16934 8881 16944 9034
rect 17050 8881 17060 9034
rect 17126 8881 17136 9034
rect 17242 8881 17252 9034
rect 17318 8881 17328 9034
rect 17434 8881 17444 9034
rect 17510 8881 17520 9034
rect 17626 8881 17636 9034
rect 17702 8881 17712 9034
rect 17818 8881 17828 9034
rect 17894 8881 17904 9034
rect 17940 8821 18160 9068
rect 18302 8881 18312 9034
rect 18378 8881 18388 9034
rect 18494 8881 18504 9034
rect 18570 8881 18580 9034
rect 18686 8881 18696 9034
rect 18762 8881 18772 9034
rect 18878 8881 18888 9034
rect 18954 8881 18964 9034
rect 19070 8881 19080 9034
rect 19146 8881 19156 9034
rect 19262 8881 19272 9034
rect 19338 8881 19348 9034
rect 19454 8881 19464 9034
rect 19530 8881 19540 9034
rect 19646 8881 19656 9034
rect 19722 8881 19732 9034
rect 19768 8821 19988 9068
rect 20130 8881 20140 9034
rect 20206 8881 20216 9034
rect 20322 8881 20332 9034
rect 20398 8881 20408 9034
rect 20514 8881 20524 9034
rect 20590 8881 20600 9034
rect 20706 8881 20716 9034
rect 20782 8881 20792 9034
rect 20898 8881 20908 9034
rect 20974 8881 20984 9034
rect 21090 8881 21100 9034
rect 21166 8881 21176 9034
rect 21282 8881 21292 9034
rect 21358 8881 21368 9034
rect 21474 8881 21484 9034
rect 21550 8881 21560 9034
rect 21596 8821 21816 9068
rect 118 8668 128 8821
rect 194 8668 204 8821
rect 310 8668 320 8821
rect 386 8668 396 8821
rect 502 8668 512 8821
rect 578 8668 588 8821
rect 694 8668 704 8821
rect 770 8668 780 8821
rect 886 8668 896 8821
rect 962 8668 972 8821
rect 1078 8668 1088 8821
rect 1154 8668 1164 8821
rect 1270 8668 1280 8821
rect 1346 8668 1356 8821
rect 1462 8668 1472 8821
rect 1528 8668 1708 8821
rect 1946 8668 1956 8821
rect 2022 8668 2032 8821
rect 2138 8668 2148 8821
rect 2214 8668 2224 8821
rect 2330 8668 2340 8821
rect 2406 8668 2416 8821
rect 2522 8668 2532 8821
rect 2598 8668 2608 8821
rect 2714 8668 2724 8821
rect 2790 8668 2800 8821
rect 2906 8668 2916 8821
rect 2982 8668 2992 8821
rect 3098 8668 3108 8821
rect 3174 8668 3184 8821
rect 3290 8668 3300 8821
rect 3356 8668 3536 8821
rect 3774 8668 3784 8821
rect 3850 8668 3860 8821
rect 3966 8668 3976 8821
rect 4042 8668 4052 8821
rect 4158 8668 4168 8821
rect 4234 8668 4244 8821
rect 4350 8668 4360 8821
rect 4426 8668 4436 8821
rect 4542 8668 4552 8821
rect 4618 8668 4628 8821
rect 4734 8668 4744 8821
rect 4810 8668 4820 8821
rect 4926 8668 4936 8821
rect 5002 8668 5012 8821
rect 5118 8668 5128 8821
rect 5184 8668 5364 8821
rect 5602 8668 5612 8821
rect 5678 8668 5688 8821
rect 5794 8668 5804 8821
rect 5870 8668 5880 8821
rect 5986 8668 5996 8821
rect 6062 8668 6072 8821
rect 6178 8668 6188 8821
rect 6254 8668 6264 8821
rect 6370 8668 6380 8821
rect 6446 8668 6456 8821
rect 6562 8668 6572 8821
rect 6638 8668 6648 8821
rect 6754 8668 6764 8821
rect 6830 8668 6840 8821
rect 6946 8668 6956 8821
rect 7012 8668 7192 8821
rect 7430 8668 7440 8821
rect 7506 8668 7516 8821
rect 7622 8668 7632 8821
rect 7698 8668 7708 8821
rect 7814 8668 7824 8821
rect 7890 8668 7900 8821
rect 8006 8668 8016 8821
rect 8082 8668 8092 8821
rect 8198 8668 8208 8821
rect 8274 8668 8284 8821
rect 8390 8668 8400 8821
rect 8466 8668 8476 8821
rect 8582 8668 8592 8821
rect 8658 8668 8668 8821
rect 8774 8668 8784 8821
rect 8840 8668 9020 8821
rect 9258 8668 9268 8821
rect 9334 8668 9344 8821
rect 9450 8668 9460 8821
rect 9526 8668 9536 8821
rect 9642 8668 9652 8821
rect 9718 8668 9728 8821
rect 9834 8668 9844 8821
rect 9910 8668 9920 8821
rect 10026 8668 10036 8821
rect 10102 8668 10112 8821
rect 10218 8668 10228 8821
rect 10294 8668 10304 8821
rect 10410 8668 10420 8821
rect 10486 8668 10496 8821
rect 10602 8668 10612 8821
rect 10668 8668 10848 8821
rect 11086 8668 11096 8821
rect 11162 8668 11172 8821
rect 11278 8668 11288 8821
rect 11354 8668 11364 8821
rect 11470 8668 11480 8821
rect 11546 8668 11556 8821
rect 11662 8668 11672 8821
rect 11738 8668 11748 8821
rect 11854 8668 11864 8821
rect 11930 8668 11940 8821
rect 12046 8668 12056 8821
rect 12122 8668 12132 8821
rect 12238 8668 12248 8821
rect 12314 8668 12324 8821
rect 12430 8668 12440 8821
rect 12496 8668 12676 8821
rect 12914 8668 12924 8821
rect 12990 8668 13000 8821
rect 13106 8668 13116 8821
rect 13182 8668 13192 8821
rect 13298 8668 13308 8821
rect 13374 8668 13384 8821
rect 13490 8668 13500 8821
rect 13566 8668 13576 8821
rect 13682 8668 13692 8821
rect 13758 8668 13768 8821
rect 13874 8668 13884 8821
rect 13950 8668 13960 8821
rect 14066 8668 14076 8821
rect 14142 8668 14152 8821
rect 14258 8668 14268 8821
rect 14324 8668 14504 8821
rect 14742 8668 14752 8821
rect 14818 8668 14828 8821
rect 14934 8668 14944 8821
rect 15010 8668 15020 8821
rect 15126 8668 15136 8821
rect 15202 8668 15212 8821
rect 15318 8668 15328 8821
rect 15394 8668 15404 8821
rect 15510 8668 15520 8821
rect 15586 8668 15596 8821
rect 15702 8668 15712 8821
rect 15778 8668 15788 8821
rect 15894 8668 15904 8821
rect 15970 8668 15980 8821
rect 16086 8668 16096 8821
rect 16152 8668 16332 8821
rect 16570 8668 16580 8821
rect 16646 8668 16656 8821
rect 16762 8668 16772 8821
rect 16838 8668 16848 8821
rect 16954 8668 16964 8821
rect 17030 8668 17040 8821
rect 17146 8668 17156 8821
rect 17222 8668 17232 8821
rect 17338 8668 17348 8821
rect 17414 8668 17424 8821
rect 17530 8668 17540 8821
rect 17606 8668 17616 8821
rect 17722 8668 17732 8821
rect 17798 8668 17808 8821
rect 17914 8668 17924 8821
rect 17980 8668 18160 8821
rect 18398 8668 18408 8821
rect 18474 8668 18484 8821
rect 18590 8668 18600 8821
rect 18666 8668 18676 8821
rect 18782 8668 18792 8821
rect 18858 8668 18868 8821
rect 18974 8668 18984 8821
rect 19050 8668 19060 8821
rect 19166 8668 19176 8821
rect 19242 8668 19252 8821
rect 19358 8668 19368 8821
rect 19434 8668 19444 8821
rect 19550 8668 19560 8821
rect 19626 8668 19636 8821
rect 19742 8668 19752 8821
rect 19808 8668 19988 8821
rect 20226 8668 20236 8821
rect 20302 8668 20312 8821
rect 20418 8668 20428 8821
rect 20494 8668 20504 8821
rect 20610 8668 20620 8821
rect 20686 8668 20696 8821
rect 20802 8668 20812 8821
rect 20878 8668 20888 8821
rect 20994 8668 21004 8821
rect 21070 8668 21080 8821
rect 21186 8668 21196 8821
rect 21262 8668 21272 8821
rect 21378 8668 21388 8821
rect 21454 8668 21464 8821
rect 21570 8668 21580 8821
rect 21636 8668 21816 8821
rect 0 8571 1490 8630
rect 1828 8571 3318 8630
rect 3656 8571 5146 8630
rect 5484 8571 6974 8630
rect 7312 8571 8802 8630
rect 9140 8571 10630 8630
rect 10968 8571 12458 8630
rect 12796 8571 14286 8630
rect 14624 8571 16114 8630
rect 16452 8571 17942 8630
rect 18280 8571 19770 8630
rect 20108 8571 21598 8630
rect 0 8392 1490 8451
rect 1828 8392 3318 8451
rect 3656 8392 5146 8451
rect 5484 8392 6974 8451
rect 7312 8392 8802 8451
rect 9140 8392 10630 8451
rect 10968 8392 12458 8451
rect 12796 8392 14286 8451
rect 14624 8392 16114 8451
rect 16452 8392 17942 8451
rect 18280 8392 19770 8451
rect 20108 8392 21598 8451
rect 22 8167 32 8320
rect 98 8167 108 8320
rect 214 8167 224 8320
rect 290 8167 300 8320
rect 406 8167 416 8320
rect 482 8167 492 8320
rect 598 8167 608 8320
rect 674 8167 684 8320
rect 790 8167 800 8320
rect 866 8167 876 8320
rect 982 8167 992 8320
rect 1058 8167 1068 8320
rect 1174 8167 1184 8320
rect 1250 8167 1260 8320
rect 1366 8167 1376 8320
rect 1442 8167 1452 8320
rect 1488 8107 1708 8354
rect 1850 8167 1860 8320
rect 1926 8167 1936 8320
rect 2042 8167 2052 8320
rect 2118 8167 2128 8320
rect 2234 8167 2244 8320
rect 2310 8167 2320 8320
rect 2426 8167 2436 8320
rect 2502 8167 2512 8320
rect 2618 8167 2628 8320
rect 2694 8167 2704 8320
rect 2810 8167 2820 8320
rect 2886 8167 2896 8320
rect 3002 8167 3012 8320
rect 3078 8167 3088 8320
rect 3194 8167 3204 8320
rect 3270 8167 3280 8320
rect 3316 8107 3536 8354
rect 3678 8167 3688 8320
rect 3754 8167 3764 8320
rect 3870 8167 3880 8320
rect 3946 8167 3956 8320
rect 4062 8167 4072 8320
rect 4138 8167 4148 8320
rect 4254 8167 4264 8320
rect 4330 8167 4340 8320
rect 4446 8167 4456 8320
rect 4522 8167 4532 8320
rect 4638 8167 4648 8320
rect 4714 8167 4724 8320
rect 4830 8167 4840 8320
rect 4906 8167 4916 8320
rect 5022 8167 5032 8320
rect 5098 8167 5108 8320
rect 5144 8107 5364 8354
rect 5506 8167 5516 8320
rect 5582 8167 5592 8320
rect 5698 8167 5708 8320
rect 5774 8167 5784 8320
rect 5890 8167 5900 8320
rect 5966 8167 5976 8320
rect 6082 8167 6092 8320
rect 6158 8167 6168 8320
rect 6274 8167 6284 8320
rect 6350 8167 6360 8320
rect 6466 8167 6476 8320
rect 6542 8167 6552 8320
rect 6658 8167 6668 8320
rect 6734 8167 6744 8320
rect 6850 8167 6860 8320
rect 6926 8167 6936 8320
rect 6972 8107 7192 8354
rect 7334 8167 7344 8320
rect 7410 8167 7420 8320
rect 7526 8167 7536 8320
rect 7602 8167 7612 8320
rect 7718 8167 7728 8320
rect 7794 8167 7804 8320
rect 7910 8167 7920 8320
rect 7986 8167 7996 8320
rect 8102 8167 8112 8320
rect 8178 8167 8188 8320
rect 8294 8167 8304 8320
rect 8370 8167 8380 8320
rect 8486 8167 8496 8320
rect 8562 8167 8572 8320
rect 8678 8167 8688 8320
rect 8754 8167 8764 8320
rect 8800 8107 9020 8354
rect 9162 8167 9172 8320
rect 9238 8167 9248 8320
rect 9354 8167 9364 8320
rect 9430 8167 9440 8320
rect 9546 8167 9556 8320
rect 9622 8167 9632 8320
rect 9738 8167 9748 8320
rect 9814 8167 9824 8320
rect 9930 8167 9940 8320
rect 10006 8167 10016 8320
rect 10122 8167 10132 8320
rect 10198 8167 10208 8320
rect 10314 8167 10324 8320
rect 10390 8167 10400 8320
rect 10506 8167 10516 8320
rect 10582 8167 10592 8320
rect 10628 8107 10848 8354
rect 10990 8167 11000 8320
rect 11066 8167 11076 8320
rect 11182 8167 11192 8320
rect 11258 8167 11268 8320
rect 11374 8167 11384 8320
rect 11450 8167 11460 8320
rect 11566 8167 11576 8320
rect 11642 8167 11652 8320
rect 11758 8167 11768 8320
rect 11834 8167 11844 8320
rect 11950 8167 11960 8320
rect 12026 8167 12036 8320
rect 12142 8167 12152 8320
rect 12218 8167 12228 8320
rect 12334 8167 12344 8320
rect 12410 8167 12420 8320
rect 12456 8107 12676 8354
rect 12818 8167 12828 8320
rect 12894 8167 12904 8320
rect 13010 8167 13020 8320
rect 13086 8167 13096 8320
rect 13202 8167 13212 8320
rect 13278 8167 13288 8320
rect 13394 8167 13404 8320
rect 13470 8167 13480 8320
rect 13586 8167 13596 8320
rect 13662 8167 13672 8320
rect 13778 8167 13788 8320
rect 13854 8167 13864 8320
rect 13970 8167 13980 8320
rect 14046 8167 14056 8320
rect 14162 8167 14172 8320
rect 14238 8167 14248 8320
rect 14284 8107 14504 8354
rect 14646 8167 14656 8320
rect 14722 8167 14732 8320
rect 14838 8167 14848 8320
rect 14914 8167 14924 8320
rect 15030 8167 15040 8320
rect 15106 8167 15116 8320
rect 15222 8167 15232 8320
rect 15298 8167 15308 8320
rect 15414 8167 15424 8320
rect 15490 8167 15500 8320
rect 15606 8167 15616 8320
rect 15682 8167 15692 8320
rect 15798 8167 15808 8320
rect 15874 8167 15884 8320
rect 15990 8167 16000 8320
rect 16066 8167 16076 8320
rect 16112 8107 16332 8354
rect 16474 8167 16484 8320
rect 16550 8167 16560 8320
rect 16666 8167 16676 8320
rect 16742 8167 16752 8320
rect 16858 8167 16868 8320
rect 16934 8167 16944 8320
rect 17050 8167 17060 8320
rect 17126 8167 17136 8320
rect 17242 8167 17252 8320
rect 17318 8167 17328 8320
rect 17434 8167 17444 8320
rect 17510 8167 17520 8320
rect 17626 8167 17636 8320
rect 17702 8167 17712 8320
rect 17818 8167 17828 8320
rect 17894 8167 17904 8320
rect 17940 8107 18160 8354
rect 18302 8167 18312 8320
rect 18378 8167 18388 8320
rect 18494 8167 18504 8320
rect 18570 8167 18580 8320
rect 18686 8167 18696 8320
rect 18762 8167 18772 8320
rect 18878 8167 18888 8320
rect 18954 8167 18964 8320
rect 19070 8167 19080 8320
rect 19146 8167 19156 8320
rect 19262 8167 19272 8320
rect 19338 8167 19348 8320
rect 19454 8167 19464 8320
rect 19530 8167 19540 8320
rect 19646 8167 19656 8320
rect 19722 8167 19732 8320
rect 19768 8107 19988 8354
rect 20130 8167 20140 8320
rect 20206 8167 20216 8320
rect 20322 8167 20332 8320
rect 20398 8167 20408 8320
rect 20514 8167 20524 8320
rect 20590 8167 20600 8320
rect 20706 8167 20716 8320
rect 20782 8167 20792 8320
rect 20898 8167 20908 8320
rect 20974 8167 20984 8320
rect 21090 8167 21100 8320
rect 21166 8167 21176 8320
rect 21282 8167 21292 8320
rect 21358 8167 21368 8320
rect 21474 8167 21484 8320
rect 21550 8167 21560 8320
rect 21596 8107 21816 8354
rect 118 7954 128 8107
rect 194 7954 204 8107
rect 310 7954 320 8107
rect 386 7954 396 8107
rect 502 7954 512 8107
rect 578 7954 588 8107
rect 694 7954 704 8107
rect 770 7954 780 8107
rect 886 7954 896 8107
rect 962 7954 972 8107
rect 1078 7954 1088 8107
rect 1154 7954 1164 8107
rect 1270 7954 1280 8107
rect 1346 7954 1356 8107
rect 1462 7954 1472 8107
rect 1528 7954 1708 8107
rect 1946 7954 1956 8107
rect 2022 7954 2032 8107
rect 2138 7954 2148 8107
rect 2214 7954 2224 8107
rect 2330 7954 2340 8107
rect 2406 7954 2416 8107
rect 2522 7954 2532 8107
rect 2598 7954 2608 8107
rect 2714 7954 2724 8107
rect 2790 7954 2800 8107
rect 2906 7954 2916 8107
rect 2982 7954 2992 8107
rect 3098 7954 3108 8107
rect 3174 7954 3184 8107
rect 3290 7954 3300 8107
rect 3356 7954 3536 8107
rect 3774 7954 3784 8107
rect 3850 7954 3860 8107
rect 3966 7954 3976 8107
rect 4042 7954 4052 8107
rect 4158 7954 4168 8107
rect 4234 7954 4244 8107
rect 4350 7954 4360 8107
rect 4426 7954 4436 8107
rect 4542 7954 4552 8107
rect 4618 7954 4628 8107
rect 4734 7954 4744 8107
rect 4810 7954 4820 8107
rect 4926 7954 4936 8107
rect 5002 7954 5012 8107
rect 5118 7954 5128 8107
rect 5184 7954 5364 8107
rect 5602 7954 5612 8107
rect 5678 7954 5688 8107
rect 5794 7954 5804 8107
rect 5870 7954 5880 8107
rect 5986 7954 5996 8107
rect 6062 7954 6072 8107
rect 6178 7954 6188 8107
rect 6254 7954 6264 8107
rect 6370 7954 6380 8107
rect 6446 7954 6456 8107
rect 6562 7954 6572 8107
rect 6638 7954 6648 8107
rect 6754 7954 6764 8107
rect 6830 7954 6840 8107
rect 6946 7954 6956 8107
rect 7012 7954 7192 8107
rect 7430 7954 7440 8107
rect 7506 7954 7516 8107
rect 7622 7954 7632 8107
rect 7698 7954 7708 8107
rect 7814 7954 7824 8107
rect 7890 7954 7900 8107
rect 8006 7954 8016 8107
rect 8082 7954 8092 8107
rect 8198 7954 8208 8107
rect 8274 7954 8284 8107
rect 8390 7954 8400 8107
rect 8466 7954 8476 8107
rect 8582 7954 8592 8107
rect 8658 7954 8668 8107
rect 8774 7954 8784 8107
rect 8840 7954 9020 8107
rect 9258 7954 9268 8107
rect 9334 7954 9344 8107
rect 9450 7954 9460 8107
rect 9526 7954 9536 8107
rect 9642 7954 9652 8107
rect 9718 7954 9728 8107
rect 9834 7954 9844 8107
rect 9910 7954 9920 8107
rect 10026 7954 10036 8107
rect 10102 7954 10112 8107
rect 10218 7954 10228 8107
rect 10294 7954 10304 8107
rect 10410 7954 10420 8107
rect 10486 7954 10496 8107
rect 10602 7954 10612 8107
rect 10668 7954 10848 8107
rect 11086 7954 11096 8107
rect 11162 7954 11172 8107
rect 11278 7954 11288 8107
rect 11354 7954 11364 8107
rect 11470 7954 11480 8107
rect 11546 7954 11556 8107
rect 11662 7954 11672 8107
rect 11738 7954 11748 8107
rect 11854 7954 11864 8107
rect 11930 7954 11940 8107
rect 12046 7954 12056 8107
rect 12122 7954 12132 8107
rect 12238 7954 12248 8107
rect 12314 7954 12324 8107
rect 12430 7954 12440 8107
rect 12496 7954 12676 8107
rect 12914 7954 12924 8107
rect 12990 7954 13000 8107
rect 13106 7954 13116 8107
rect 13182 7954 13192 8107
rect 13298 7954 13308 8107
rect 13374 7954 13384 8107
rect 13490 7954 13500 8107
rect 13566 7954 13576 8107
rect 13682 7954 13692 8107
rect 13758 7954 13768 8107
rect 13874 7954 13884 8107
rect 13950 7954 13960 8107
rect 14066 7954 14076 8107
rect 14142 7954 14152 8107
rect 14258 7954 14268 8107
rect 14324 7954 14504 8107
rect 14742 7954 14752 8107
rect 14818 7954 14828 8107
rect 14934 7954 14944 8107
rect 15010 7954 15020 8107
rect 15126 7954 15136 8107
rect 15202 7954 15212 8107
rect 15318 7954 15328 8107
rect 15394 7954 15404 8107
rect 15510 7954 15520 8107
rect 15586 7954 15596 8107
rect 15702 7954 15712 8107
rect 15778 7954 15788 8107
rect 15894 7954 15904 8107
rect 15970 7954 15980 8107
rect 16086 7954 16096 8107
rect 16152 7954 16332 8107
rect 16570 7954 16580 8107
rect 16646 7954 16656 8107
rect 16762 7954 16772 8107
rect 16838 7954 16848 8107
rect 16954 7954 16964 8107
rect 17030 7954 17040 8107
rect 17146 7954 17156 8107
rect 17222 7954 17232 8107
rect 17338 7954 17348 8107
rect 17414 7954 17424 8107
rect 17530 7954 17540 8107
rect 17606 7954 17616 8107
rect 17722 7954 17732 8107
rect 17798 7954 17808 8107
rect 17914 7954 17924 8107
rect 17980 7954 18160 8107
rect 18398 7954 18408 8107
rect 18474 7954 18484 8107
rect 18590 7954 18600 8107
rect 18666 7954 18676 8107
rect 18782 7954 18792 8107
rect 18858 7954 18868 8107
rect 18974 7954 18984 8107
rect 19050 7954 19060 8107
rect 19166 7954 19176 8107
rect 19242 7954 19252 8107
rect 19358 7954 19368 8107
rect 19434 7954 19444 8107
rect 19550 7954 19560 8107
rect 19626 7954 19636 8107
rect 19742 7954 19752 8107
rect 19808 7954 19988 8107
rect 20226 7954 20236 8107
rect 20302 7954 20312 8107
rect 20418 7954 20428 8107
rect 20494 7954 20504 8107
rect 20610 7954 20620 8107
rect 20686 7954 20696 8107
rect 20802 7954 20812 8107
rect 20878 7954 20888 8107
rect 20994 7954 21004 8107
rect 21070 7954 21080 8107
rect 21186 7954 21196 8107
rect 21262 7954 21272 8107
rect 21378 7954 21388 8107
rect 21454 7954 21464 8107
rect 21570 7954 21580 8107
rect 21636 7954 21816 8107
rect 0 7857 1490 7916
rect 1828 7857 3318 7916
rect 3656 7857 5146 7916
rect 5484 7857 6974 7916
rect 7312 7857 8802 7916
rect 9140 7857 10630 7916
rect 10968 7857 12458 7916
rect 12796 7857 14286 7916
rect 14624 7857 16114 7916
rect 16452 7857 17942 7916
rect 18280 7857 19770 7916
rect 20108 7857 21598 7916
rect 0 7678 1490 7737
rect 1828 7678 3318 7737
rect 3656 7678 5146 7737
rect 5484 7678 6974 7737
rect 7312 7678 8802 7737
rect 9140 7678 10630 7737
rect 10968 7678 12458 7737
rect 12796 7678 14286 7737
rect 14624 7678 16114 7737
rect 16452 7678 17942 7737
rect 18280 7678 19770 7737
rect 20108 7678 21598 7737
rect 22 7453 32 7606
rect 98 7453 108 7606
rect 214 7453 224 7606
rect 290 7453 300 7606
rect 406 7453 416 7606
rect 482 7453 492 7606
rect 598 7453 608 7606
rect 674 7453 684 7606
rect 790 7453 800 7606
rect 866 7453 876 7606
rect 982 7453 992 7606
rect 1058 7453 1068 7606
rect 1174 7453 1184 7606
rect 1250 7453 1260 7606
rect 1366 7453 1376 7606
rect 1442 7453 1452 7606
rect 1488 7393 1708 7640
rect 1850 7453 1860 7606
rect 1926 7453 1936 7606
rect 2042 7453 2052 7606
rect 2118 7453 2128 7606
rect 2234 7453 2244 7606
rect 2310 7453 2320 7606
rect 2426 7453 2436 7606
rect 2502 7453 2512 7606
rect 2618 7453 2628 7606
rect 2694 7453 2704 7606
rect 2810 7453 2820 7606
rect 2886 7453 2896 7606
rect 3002 7453 3012 7606
rect 3078 7453 3088 7606
rect 3194 7453 3204 7606
rect 3270 7453 3280 7606
rect 3316 7393 3536 7640
rect 3678 7453 3688 7606
rect 3754 7453 3764 7606
rect 3870 7453 3880 7606
rect 3946 7453 3956 7606
rect 4062 7453 4072 7606
rect 4138 7453 4148 7606
rect 4254 7453 4264 7606
rect 4330 7453 4340 7606
rect 4446 7453 4456 7606
rect 4522 7453 4532 7606
rect 4638 7453 4648 7606
rect 4714 7453 4724 7606
rect 4830 7453 4840 7606
rect 4906 7453 4916 7606
rect 5022 7453 5032 7606
rect 5098 7453 5108 7606
rect 5144 7393 5364 7640
rect 5506 7453 5516 7606
rect 5582 7453 5592 7606
rect 5698 7453 5708 7606
rect 5774 7453 5784 7606
rect 5890 7453 5900 7606
rect 5966 7453 5976 7606
rect 6082 7453 6092 7606
rect 6158 7453 6168 7606
rect 6274 7453 6284 7606
rect 6350 7453 6360 7606
rect 6466 7453 6476 7606
rect 6542 7453 6552 7606
rect 6658 7453 6668 7606
rect 6734 7453 6744 7606
rect 6850 7453 6860 7606
rect 6926 7453 6936 7606
rect 6972 7393 7192 7640
rect 7334 7453 7344 7606
rect 7410 7453 7420 7606
rect 7526 7453 7536 7606
rect 7602 7453 7612 7606
rect 7718 7453 7728 7606
rect 7794 7453 7804 7606
rect 7910 7453 7920 7606
rect 7986 7453 7996 7606
rect 8102 7453 8112 7606
rect 8178 7453 8188 7606
rect 8294 7453 8304 7606
rect 8370 7453 8380 7606
rect 8486 7453 8496 7606
rect 8562 7453 8572 7606
rect 8678 7453 8688 7606
rect 8754 7453 8764 7606
rect 8800 7393 9020 7640
rect 9162 7453 9172 7606
rect 9238 7453 9248 7606
rect 9354 7453 9364 7606
rect 9430 7453 9440 7606
rect 9546 7453 9556 7606
rect 9622 7453 9632 7606
rect 9738 7453 9748 7606
rect 9814 7453 9824 7606
rect 9930 7453 9940 7606
rect 10006 7453 10016 7606
rect 10122 7453 10132 7606
rect 10198 7453 10208 7606
rect 10314 7453 10324 7606
rect 10390 7453 10400 7606
rect 10506 7453 10516 7606
rect 10582 7453 10592 7606
rect 10628 7393 10848 7640
rect 10990 7453 11000 7606
rect 11066 7453 11076 7606
rect 11182 7453 11192 7606
rect 11258 7453 11268 7606
rect 11374 7453 11384 7606
rect 11450 7453 11460 7606
rect 11566 7453 11576 7606
rect 11642 7453 11652 7606
rect 11758 7453 11768 7606
rect 11834 7453 11844 7606
rect 11950 7453 11960 7606
rect 12026 7453 12036 7606
rect 12142 7453 12152 7606
rect 12218 7453 12228 7606
rect 12334 7453 12344 7606
rect 12410 7453 12420 7606
rect 12456 7393 12676 7640
rect 12818 7453 12828 7606
rect 12894 7453 12904 7606
rect 13010 7453 13020 7606
rect 13086 7453 13096 7606
rect 13202 7453 13212 7606
rect 13278 7453 13288 7606
rect 13394 7453 13404 7606
rect 13470 7453 13480 7606
rect 13586 7453 13596 7606
rect 13662 7453 13672 7606
rect 13778 7453 13788 7606
rect 13854 7453 13864 7606
rect 13970 7453 13980 7606
rect 14046 7453 14056 7606
rect 14162 7453 14172 7606
rect 14238 7453 14248 7606
rect 14284 7393 14504 7640
rect 14646 7453 14656 7606
rect 14722 7453 14732 7606
rect 14838 7453 14848 7606
rect 14914 7453 14924 7606
rect 15030 7453 15040 7606
rect 15106 7453 15116 7606
rect 15222 7453 15232 7606
rect 15298 7453 15308 7606
rect 15414 7453 15424 7606
rect 15490 7453 15500 7606
rect 15606 7453 15616 7606
rect 15682 7453 15692 7606
rect 15798 7453 15808 7606
rect 15874 7453 15884 7606
rect 15990 7453 16000 7606
rect 16066 7453 16076 7606
rect 16112 7393 16332 7640
rect 16474 7453 16484 7606
rect 16550 7453 16560 7606
rect 16666 7453 16676 7606
rect 16742 7453 16752 7606
rect 16858 7453 16868 7606
rect 16934 7453 16944 7606
rect 17050 7453 17060 7606
rect 17126 7453 17136 7606
rect 17242 7453 17252 7606
rect 17318 7453 17328 7606
rect 17434 7453 17444 7606
rect 17510 7453 17520 7606
rect 17626 7453 17636 7606
rect 17702 7453 17712 7606
rect 17818 7453 17828 7606
rect 17894 7453 17904 7606
rect 17940 7393 18160 7640
rect 18302 7453 18312 7606
rect 18378 7453 18388 7606
rect 18494 7453 18504 7606
rect 18570 7453 18580 7606
rect 18686 7453 18696 7606
rect 18762 7453 18772 7606
rect 18878 7453 18888 7606
rect 18954 7453 18964 7606
rect 19070 7453 19080 7606
rect 19146 7453 19156 7606
rect 19262 7453 19272 7606
rect 19338 7453 19348 7606
rect 19454 7453 19464 7606
rect 19530 7453 19540 7606
rect 19646 7453 19656 7606
rect 19722 7453 19732 7606
rect 19768 7393 19988 7640
rect 20130 7453 20140 7606
rect 20206 7453 20216 7606
rect 20322 7453 20332 7606
rect 20398 7453 20408 7606
rect 20514 7453 20524 7606
rect 20590 7453 20600 7606
rect 20706 7453 20716 7606
rect 20782 7453 20792 7606
rect 20898 7453 20908 7606
rect 20974 7453 20984 7606
rect 21090 7453 21100 7606
rect 21166 7453 21176 7606
rect 21282 7453 21292 7606
rect 21358 7453 21368 7606
rect 21474 7453 21484 7606
rect 21550 7453 21560 7606
rect 21596 7393 21816 7640
rect 118 7240 128 7393
rect 194 7240 204 7393
rect 310 7240 320 7393
rect 386 7240 396 7393
rect 502 7240 512 7393
rect 578 7240 588 7393
rect 694 7240 704 7393
rect 770 7240 780 7393
rect 886 7240 896 7393
rect 962 7240 972 7393
rect 1078 7240 1088 7393
rect 1154 7240 1164 7393
rect 1270 7240 1280 7393
rect 1346 7240 1356 7393
rect 1462 7240 1472 7393
rect 1528 7240 1708 7393
rect 1946 7240 1956 7393
rect 2022 7240 2032 7393
rect 2138 7240 2148 7393
rect 2214 7240 2224 7393
rect 2330 7240 2340 7393
rect 2406 7240 2416 7393
rect 2522 7240 2532 7393
rect 2598 7240 2608 7393
rect 2714 7240 2724 7393
rect 2790 7240 2800 7393
rect 2906 7240 2916 7393
rect 2982 7240 2992 7393
rect 3098 7240 3108 7393
rect 3174 7240 3184 7393
rect 3290 7240 3300 7393
rect 3356 7240 3536 7393
rect 3774 7240 3784 7393
rect 3850 7240 3860 7393
rect 3966 7240 3976 7393
rect 4042 7240 4052 7393
rect 4158 7240 4168 7393
rect 4234 7240 4244 7393
rect 4350 7240 4360 7393
rect 4426 7240 4436 7393
rect 4542 7240 4552 7393
rect 4618 7240 4628 7393
rect 4734 7240 4744 7393
rect 4810 7240 4820 7393
rect 4926 7240 4936 7393
rect 5002 7240 5012 7393
rect 5118 7240 5128 7393
rect 5184 7240 5364 7393
rect 5602 7240 5612 7393
rect 5678 7240 5688 7393
rect 5794 7240 5804 7393
rect 5870 7240 5880 7393
rect 5986 7240 5996 7393
rect 6062 7240 6072 7393
rect 6178 7240 6188 7393
rect 6254 7240 6264 7393
rect 6370 7240 6380 7393
rect 6446 7240 6456 7393
rect 6562 7240 6572 7393
rect 6638 7240 6648 7393
rect 6754 7240 6764 7393
rect 6830 7240 6840 7393
rect 6946 7240 6956 7393
rect 7012 7240 7192 7393
rect 7430 7240 7440 7393
rect 7506 7240 7516 7393
rect 7622 7240 7632 7393
rect 7698 7240 7708 7393
rect 7814 7240 7824 7393
rect 7890 7240 7900 7393
rect 8006 7240 8016 7393
rect 8082 7240 8092 7393
rect 8198 7240 8208 7393
rect 8274 7240 8284 7393
rect 8390 7240 8400 7393
rect 8466 7240 8476 7393
rect 8582 7240 8592 7393
rect 8658 7240 8668 7393
rect 8774 7240 8784 7393
rect 8840 7240 9020 7393
rect 9258 7240 9268 7393
rect 9334 7240 9344 7393
rect 9450 7240 9460 7393
rect 9526 7240 9536 7393
rect 9642 7240 9652 7393
rect 9718 7240 9728 7393
rect 9834 7240 9844 7393
rect 9910 7240 9920 7393
rect 10026 7240 10036 7393
rect 10102 7240 10112 7393
rect 10218 7240 10228 7393
rect 10294 7240 10304 7393
rect 10410 7240 10420 7393
rect 10486 7240 10496 7393
rect 10602 7240 10612 7393
rect 10668 7240 10848 7393
rect 11086 7240 11096 7393
rect 11162 7240 11172 7393
rect 11278 7240 11288 7393
rect 11354 7240 11364 7393
rect 11470 7240 11480 7393
rect 11546 7240 11556 7393
rect 11662 7240 11672 7393
rect 11738 7240 11748 7393
rect 11854 7240 11864 7393
rect 11930 7240 11940 7393
rect 12046 7240 12056 7393
rect 12122 7240 12132 7393
rect 12238 7240 12248 7393
rect 12314 7240 12324 7393
rect 12430 7240 12440 7393
rect 12496 7240 12676 7393
rect 12914 7240 12924 7393
rect 12990 7240 13000 7393
rect 13106 7240 13116 7393
rect 13182 7240 13192 7393
rect 13298 7240 13308 7393
rect 13374 7240 13384 7393
rect 13490 7240 13500 7393
rect 13566 7240 13576 7393
rect 13682 7240 13692 7393
rect 13758 7240 13768 7393
rect 13874 7240 13884 7393
rect 13950 7240 13960 7393
rect 14066 7240 14076 7393
rect 14142 7240 14152 7393
rect 14258 7240 14268 7393
rect 14324 7240 14504 7393
rect 14742 7240 14752 7393
rect 14818 7240 14828 7393
rect 14934 7240 14944 7393
rect 15010 7240 15020 7393
rect 15126 7240 15136 7393
rect 15202 7240 15212 7393
rect 15318 7240 15328 7393
rect 15394 7240 15404 7393
rect 15510 7240 15520 7393
rect 15586 7240 15596 7393
rect 15702 7240 15712 7393
rect 15778 7240 15788 7393
rect 15894 7240 15904 7393
rect 15970 7240 15980 7393
rect 16086 7240 16096 7393
rect 16152 7240 16332 7393
rect 16570 7240 16580 7393
rect 16646 7240 16656 7393
rect 16762 7240 16772 7393
rect 16838 7240 16848 7393
rect 16954 7240 16964 7393
rect 17030 7240 17040 7393
rect 17146 7240 17156 7393
rect 17222 7240 17232 7393
rect 17338 7240 17348 7393
rect 17414 7240 17424 7393
rect 17530 7240 17540 7393
rect 17606 7240 17616 7393
rect 17722 7240 17732 7393
rect 17798 7240 17808 7393
rect 17914 7240 17924 7393
rect 17980 7240 18160 7393
rect 18398 7240 18408 7393
rect 18474 7240 18484 7393
rect 18590 7240 18600 7393
rect 18666 7240 18676 7393
rect 18782 7240 18792 7393
rect 18858 7240 18868 7393
rect 18974 7240 18984 7393
rect 19050 7240 19060 7393
rect 19166 7240 19176 7393
rect 19242 7240 19252 7393
rect 19358 7240 19368 7393
rect 19434 7240 19444 7393
rect 19550 7240 19560 7393
rect 19626 7240 19636 7393
rect 19742 7240 19752 7393
rect 19808 7240 19988 7393
rect 20226 7240 20236 7393
rect 20302 7240 20312 7393
rect 20418 7240 20428 7393
rect 20494 7240 20504 7393
rect 20610 7240 20620 7393
rect 20686 7240 20696 7393
rect 20802 7240 20812 7393
rect 20878 7240 20888 7393
rect 20994 7240 21004 7393
rect 21070 7240 21080 7393
rect 21186 7240 21196 7393
rect 21262 7240 21272 7393
rect 21378 7240 21388 7393
rect 21454 7240 21464 7393
rect 21570 7240 21580 7393
rect 21636 7240 21816 7393
rect 0 7143 1490 7202
rect 1828 7143 3318 7202
rect 3656 7143 5146 7202
rect 5484 7143 6974 7202
rect 7312 7143 8802 7202
rect 9140 7143 10630 7202
rect 10968 7143 12458 7202
rect 12796 7143 14286 7202
rect 14624 7143 16114 7202
rect 16452 7143 17942 7202
rect 18280 7143 19770 7202
rect 20108 7143 21598 7202
rect 0 6964 1490 7023
rect 1828 6964 3318 7023
rect 3656 6964 5146 7023
rect 5484 6964 6974 7023
rect 7312 6964 8802 7023
rect 9140 6964 10630 7023
rect 10968 6964 12458 7023
rect 12796 6964 14286 7023
rect 14624 6964 16114 7023
rect 16452 6964 17942 7023
rect 18280 6964 19770 7023
rect 20108 6964 21598 7023
rect 22 6739 32 6892
rect 98 6739 108 6892
rect 214 6739 224 6892
rect 290 6739 300 6892
rect 406 6739 416 6892
rect 482 6739 492 6892
rect 598 6739 608 6892
rect 674 6739 684 6892
rect 790 6739 800 6892
rect 866 6739 876 6892
rect 982 6739 992 6892
rect 1058 6739 1068 6892
rect 1174 6739 1184 6892
rect 1250 6739 1260 6892
rect 1366 6739 1376 6892
rect 1442 6739 1452 6892
rect 1488 6679 1708 6926
rect 1850 6739 1860 6892
rect 1926 6739 1936 6892
rect 2042 6739 2052 6892
rect 2118 6739 2128 6892
rect 2234 6739 2244 6892
rect 2310 6739 2320 6892
rect 2426 6739 2436 6892
rect 2502 6739 2512 6892
rect 2618 6739 2628 6892
rect 2694 6739 2704 6892
rect 2810 6739 2820 6892
rect 2886 6739 2896 6892
rect 3002 6739 3012 6892
rect 3078 6739 3088 6892
rect 3194 6739 3204 6892
rect 3270 6739 3280 6892
rect 3316 6679 3536 6926
rect 3678 6739 3688 6892
rect 3754 6739 3764 6892
rect 3870 6739 3880 6892
rect 3946 6739 3956 6892
rect 4062 6739 4072 6892
rect 4138 6739 4148 6892
rect 4254 6739 4264 6892
rect 4330 6739 4340 6892
rect 4446 6739 4456 6892
rect 4522 6739 4532 6892
rect 4638 6739 4648 6892
rect 4714 6739 4724 6892
rect 4830 6739 4840 6892
rect 4906 6739 4916 6892
rect 5022 6739 5032 6892
rect 5098 6739 5108 6892
rect 5144 6679 5364 6926
rect 5506 6739 5516 6892
rect 5582 6739 5592 6892
rect 5698 6739 5708 6892
rect 5774 6739 5784 6892
rect 5890 6739 5900 6892
rect 5966 6739 5976 6892
rect 6082 6739 6092 6892
rect 6158 6739 6168 6892
rect 6274 6739 6284 6892
rect 6350 6739 6360 6892
rect 6466 6739 6476 6892
rect 6542 6739 6552 6892
rect 6658 6739 6668 6892
rect 6734 6739 6744 6892
rect 6850 6739 6860 6892
rect 6926 6739 6936 6892
rect 6972 6679 7192 6926
rect 7334 6739 7344 6892
rect 7410 6739 7420 6892
rect 7526 6739 7536 6892
rect 7602 6739 7612 6892
rect 7718 6739 7728 6892
rect 7794 6739 7804 6892
rect 7910 6739 7920 6892
rect 7986 6739 7996 6892
rect 8102 6739 8112 6892
rect 8178 6739 8188 6892
rect 8294 6739 8304 6892
rect 8370 6739 8380 6892
rect 8486 6739 8496 6892
rect 8562 6739 8572 6892
rect 8678 6739 8688 6892
rect 8754 6739 8764 6892
rect 8800 6679 9020 6926
rect 9162 6739 9172 6892
rect 9238 6739 9248 6892
rect 9354 6739 9364 6892
rect 9430 6739 9440 6892
rect 9546 6739 9556 6892
rect 9622 6739 9632 6892
rect 9738 6739 9748 6892
rect 9814 6739 9824 6892
rect 9930 6739 9940 6892
rect 10006 6739 10016 6892
rect 10122 6739 10132 6892
rect 10198 6739 10208 6892
rect 10314 6739 10324 6892
rect 10390 6739 10400 6892
rect 10506 6739 10516 6892
rect 10582 6739 10592 6892
rect 10628 6679 10848 6926
rect 10990 6739 11000 6892
rect 11066 6739 11076 6892
rect 11182 6739 11192 6892
rect 11258 6739 11268 6892
rect 11374 6739 11384 6892
rect 11450 6739 11460 6892
rect 11566 6739 11576 6892
rect 11642 6739 11652 6892
rect 11758 6739 11768 6892
rect 11834 6739 11844 6892
rect 11950 6739 11960 6892
rect 12026 6739 12036 6892
rect 12142 6739 12152 6892
rect 12218 6739 12228 6892
rect 12334 6739 12344 6892
rect 12410 6739 12420 6892
rect 12456 6679 12676 6926
rect 12818 6739 12828 6892
rect 12894 6739 12904 6892
rect 13010 6739 13020 6892
rect 13086 6739 13096 6892
rect 13202 6739 13212 6892
rect 13278 6739 13288 6892
rect 13394 6739 13404 6892
rect 13470 6739 13480 6892
rect 13586 6739 13596 6892
rect 13662 6739 13672 6892
rect 13778 6739 13788 6892
rect 13854 6739 13864 6892
rect 13970 6739 13980 6892
rect 14046 6739 14056 6892
rect 14162 6739 14172 6892
rect 14238 6739 14248 6892
rect 14284 6679 14504 6926
rect 14646 6739 14656 6892
rect 14722 6739 14732 6892
rect 14838 6739 14848 6892
rect 14914 6739 14924 6892
rect 15030 6739 15040 6892
rect 15106 6739 15116 6892
rect 15222 6739 15232 6892
rect 15298 6739 15308 6892
rect 15414 6739 15424 6892
rect 15490 6739 15500 6892
rect 15606 6739 15616 6892
rect 15682 6739 15692 6892
rect 15798 6739 15808 6892
rect 15874 6739 15884 6892
rect 15990 6739 16000 6892
rect 16066 6739 16076 6892
rect 16112 6679 16332 6926
rect 16474 6739 16484 6892
rect 16550 6739 16560 6892
rect 16666 6739 16676 6892
rect 16742 6739 16752 6892
rect 16858 6739 16868 6892
rect 16934 6739 16944 6892
rect 17050 6739 17060 6892
rect 17126 6739 17136 6892
rect 17242 6739 17252 6892
rect 17318 6739 17328 6892
rect 17434 6739 17444 6892
rect 17510 6739 17520 6892
rect 17626 6739 17636 6892
rect 17702 6739 17712 6892
rect 17818 6739 17828 6892
rect 17894 6739 17904 6892
rect 17940 6679 18160 6926
rect 18302 6739 18312 6892
rect 18378 6739 18388 6892
rect 18494 6739 18504 6892
rect 18570 6739 18580 6892
rect 18686 6739 18696 6892
rect 18762 6739 18772 6892
rect 18878 6739 18888 6892
rect 18954 6739 18964 6892
rect 19070 6739 19080 6892
rect 19146 6739 19156 6892
rect 19262 6739 19272 6892
rect 19338 6739 19348 6892
rect 19454 6739 19464 6892
rect 19530 6739 19540 6892
rect 19646 6739 19656 6892
rect 19722 6739 19732 6892
rect 19768 6679 19988 6926
rect 20130 6739 20140 6892
rect 20206 6739 20216 6892
rect 20322 6739 20332 6892
rect 20398 6739 20408 6892
rect 20514 6739 20524 6892
rect 20590 6739 20600 6892
rect 20706 6739 20716 6892
rect 20782 6739 20792 6892
rect 20898 6739 20908 6892
rect 20974 6739 20984 6892
rect 21090 6739 21100 6892
rect 21166 6739 21176 6892
rect 21282 6739 21292 6892
rect 21358 6739 21368 6892
rect 21474 6739 21484 6892
rect 21550 6739 21560 6892
rect 21596 6679 21816 6926
rect 118 6526 128 6679
rect 194 6526 204 6679
rect 310 6526 320 6679
rect 386 6526 396 6679
rect 502 6526 512 6679
rect 578 6526 588 6679
rect 694 6526 704 6679
rect 770 6526 780 6679
rect 886 6526 896 6679
rect 962 6526 972 6679
rect 1078 6526 1088 6679
rect 1154 6526 1164 6679
rect 1270 6526 1280 6679
rect 1346 6526 1356 6679
rect 1462 6526 1472 6679
rect 1528 6526 1708 6679
rect 1946 6526 1956 6679
rect 2022 6526 2032 6679
rect 2138 6526 2148 6679
rect 2214 6526 2224 6679
rect 2330 6526 2340 6679
rect 2406 6526 2416 6679
rect 2522 6526 2532 6679
rect 2598 6526 2608 6679
rect 2714 6526 2724 6679
rect 2790 6526 2800 6679
rect 2906 6526 2916 6679
rect 2982 6526 2992 6679
rect 3098 6526 3108 6679
rect 3174 6526 3184 6679
rect 3290 6526 3300 6679
rect 3356 6526 3536 6679
rect 3774 6526 3784 6679
rect 3850 6526 3860 6679
rect 3966 6526 3976 6679
rect 4042 6526 4052 6679
rect 4158 6526 4168 6679
rect 4234 6526 4244 6679
rect 4350 6526 4360 6679
rect 4426 6526 4436 6679
rect 4542 6526 4552 6679
rect 4618 6526 4628 6679
rect 4734 6526 4744 6679
rect 4810 6526 4820 6679
rect 4926 6526 4936 6679
rect 5002 6526 5012 6679
rect 5118 6526 5128 6679
rect 5184 6526 5364 6679
rect 5602 6526 5612 6679
rect 5678 6526 5688 6679
rect 5794 6526 5804 6679
rect 5870 6526 5880 6679
rect 5986 6526 5996 6679
rect 6062 6526 6072 6679
rect 6178 6526 6188 6679
rect 6254 6526 6264 6679
rect 6370 6526 6380 6679
rect 6446 6526 6456 6679
rect 6562 6526 6572 6679
rect 6638 6526 6648 6679
rect 6754 6526 6764 6679
rect 6830 6526 6840 6679
rect 6946 6526 6956 6679
rect 7012 6526 7192 6679
rect 7430 6526 7440 6679
rect 7506 6526 7516 6679
rect 7622 6526 7632 6679
rect 7698 6526 7708 6679
rect 7814 6526 7824 6679
rect 7890 6526 7900 6679
rect 8006 6526 8016 6679
rect 8082 6526 8092 6679
rect 8198 6526 8208 6679
rect 8274 6526 8284 6679
rect 8390 6526 8400 6679
rect 8466 6526 8476 6679
rect 8582 6526 8592 6679
rect 8658 6526 8668 6679
rect 8774 6526 8784 6679
rect 8840 6526 9020 6679
rect 9258 6526 9268 6679
rect 9334 6526 9344 6679
rect 9450 6526 9460 6679
rect 9526 6526 9536 6679
rect 9642 6526 9652 6679
rect 9718 6526 9728 6679
rect 9834 6526 9844 6679
rect 9910 6526 9920 6679
rect 10026 6526 10036 6679
rect 10102 6526 10112 6679
rect 10218 6526 10228 6679
rect 10294 6526 10304 6679
rect 10410 6526 10420 6679
rect 10486 6526 10496 6679
rect 10602 6526 10612 6679
rect 10668 6526 10848 6679
rect 11086 6526 11096 6679
rect 11162 6526 11172 6679
rect 11278 6526 11288 6679
rect 11354 6526 11364 6679
rect 11470 6526 11480 6679
rect 11546 6526 11556 6679
rect 11662 6526 11672 6679
rect 11738 6526 11748 6679
rect 11854 6526 11864 6679
rect 11930 6526 11940 6679
rect 12046 6526 12056 6679
rect 12122 6526 12132 6679
rect 12238 6526 12248 6679
rect 12314 6526 12324 6679
rect 12430 6526 12440 6679
rect 12496 6526 12676 6679
rect 12914 6526 12924 6679
rect 12990 6526 13000 6679
rect 13106 6526 13116 6679
rect 13182 6526 13192 6679
rect 13298 6526 13308 6679
rect 13374 6526 13384 6679
rect 13490 6526 13500 6679
rect 13566 6526 13576 6679
rect 13682 6526 13692 6679
rect 13758 6526 13768 6679
rect 13874 6526 13884 6679
rect 13950 6526 13960 6679
rect 14066 6526 14076 6679
rect 14142 6526 14152 6679
rect 14258 6526 14268 6679
rect 14324 6526 14504 6679
rect 14742 6526 14752 6679
rect 14818 6526 14828 6679
rect 14934 6526 14944 6679
rect 15010 6526 15020 6679
rect 15126 6526 15136 6679
rect 15202 6526 15212 6679
rect 15318 6526 15328 6679
rect 15394 6526 15404 6679
rect 15510 6526 15520 6679
rect 15586 6526 15596 6679
rect 15702 6526 15712 6679
rect 15778 6526 15788 6679
rect 15894 6526 15904 6679
rect 15970 6526 15980 6679
rect 16086 6526 16096 6679
rect 16152 6526 16332 6679
rect 16570 6526 16580 6679
rect 16646 6526 16656 6679
rect 16762 6526 16772 6679
rect 16838 6526 16848 6679
rect 16954 6526 16964 6679
rect 17030 6526 17040 6679
rect 17146 6526 17156 6679
rect 17222 6526 17232 6679
rect 17338 6526 17348 6679
rect 17414 6526 17424 6679
rect 17530 6526 17540 6679
rect 17606 6526 17616 6679
rect 17722 6526 17732 6679
rect 17798 6526 17808 6679
rect 17914 6526 17924 6679
rect 17980 6526 18160 6679
rect 18398 6526 18408 6679
rect 18474 6526 18484 6679
rect 18590 6526 18600 6679
rect 18666 6526 18676 6679
rect 18782 6526 18792 6679
rect 18858 6526 18868 6679
rect 18974 6526 18984 6679
rect 19050 6526 19060 6679
rect 19166 6526 19176 6679
rect 19242 6526 19252 6679
rect 19358 6526 19368 6679
rect 19434 6526 19444 6679
rect 19550 6526 19560 6679
rect 19626 6526 19636 6679
rect 19742 6526 19752 6679
rect 19808 6526 19988 6679
rect 20226 6526 20236 6679
rect 20302 6526 20312 6679
rect 20418 6526 20428 6679
rect 20494 6526 20504 6679
rect 20610 6526 20620 6679
rect 20686 6526 20696 6679
rect 20802 6526 20812 6679
rect 20878 6526 20888 6679
rect 20994 6526 21004 6679
rect 21070 6526 21080 6679
rect 21186 6526 21196 6679
rect 21262 6526 21272 6679
rect 21378 6526 21388 6679
rect 21454 6526 21464 6679
rect 21570 6526 21580 6679
rect 21636 6526 21816 6679
rect 0 6429 1490 6488
rect 1828 6429 3318 6488
rect 3656 6429 5146 6488
rect 5484 6429 6974 6488
rect 7312 6429 8802 6488
rect 9140 6429 10630 6488
rect 10968 6429 12458 6488
rect 12796 6429 14286 6488
rect 14624 6429 16114 6488
rect 16452 6429 17942 6488
rect 18280 6429 19770 6488
rect 20108 6429 21598 6488
rect 0 6250 1490 6309
rect 1828 6250 3318 6309
rect 3656 6250 5146 6309
rect 5484 6250 6974 6309
rect 7312 6250 8802 6309
rect 9140 6250 10630 6309
rect 10968 6250 12458 6309
rect 12796 6250 14286 6309
rect 14624 6250 16114 6309
rect 16452 6250 17942 6309
rect 18280 6250 19770 6309
rect 20108 6250 21598 6309
rect 22 6025 32 6178
rect 98 6025 108 6178
rect 214 6025 224 6178
rect 290 6025 300 6178
rect 406 6025 416 6178
rect 482 6025 492 6178
rect 598 6025 608 6178
rect 674 6025 684 6178
rect 790 6025 800 6178
rect 866 6025 876 6178
rect 982 6025 992 6178
rect 1058 6025 1068 6178
rect 1174 6025 1184 6178
rect 1250 6025 1260 6178
rect 1366 6025 1376 6178
rect 1442 6025 1452 6178
rect 1488 5965 1708 6212
rect 1850 6025 1860 6178
rect 1926 6025 1936 6178
rect 2042 6025 2052 6178
rect 2118 6025 2128 6178
rect 2234 6025 2244 6178
rect 2310 6025 2320 6178
rect 2426 6025 2436 6178
rect 2502 6025 2512 6178
rect 2618 6025 2628 6178
rect 2694 6025 2704 6178
rect 2810 6025 2820 6178
rect 2886 6025 2896 6178
rect 3002 6025 3012 6178
rect 3078 6025 3088 6178
rect 3194 6025 3204 6178
rect 3270 6025 3280 6178
rect 3316 5965 3536 6212
rect 3678 6025 3688 6178
rect 3754 6025 3764 6178
rect 3870 6025 3880 6178
rect 3946 6025 3956 6178
rect 4062 6025 4072 6178
rect 4138 6025 4148 6178
rect 4254 6025 4264 6178
rect 4330 6025 4340 6178
rect 4446 6025 4456 6178
rect 4522 6025 4532 6178
rect 4638 6025 4648 6178
rect 4714 6025 4724 6178
rect 4830 6025 4840 6178
rect 4906 6025 4916 6178
rect 5022 6025 5032 6178
rect 5098 6025 5108 6178
rect 5144 5965 5364 6212
rect 5506 6025 5516 6178
rect 5582 6025 5592 6178
rect 5698 6025 5708 6178
rect 5774 6025 5784 6178
rect 5890 6025 5900 6178
rect 5966 6025 5976 6178
rect 6082 6025 6092 6178
rect 6158 6025 6168 6178
rect 6274 6025 6284 6178
rect 6350 6025 6360 6178
rect 6466 6025 6476 6178
rect 6542 6025 6552 6178
rect 6658 6025 6668 6178
rect 6734 6025 6744 6178
rect 6850 6025 6860 6178
rect 6926 6025 6936 6178
rect 6972 5965 7192 6212
rect 7334 6025 7344 6178
rect 7410 6025 7420 6178
rect 7526 6025 7536 6178
rect 7602 6025 7612 6178
rect 7718 6025 7728 6178
rect 7794 6025 7804 6178
rect 7910 6025 7920 6178
rect 7986 6025 7996 6178
rect 8102 6025 8112 6178
rect 8178 6025 8188 6178
rect 8294 6025 8304 6178
rect 8370 6025 8380 6178
rect 8486 6025 8496 6178
rect 8562 6025 8572 6178
rect 8678 6025 8688 6178
rect 8754 6025 8764 6178
rect 8800 5965 9020 6212
rect 9162 6025 9172 6178
rect 9238 6025 9248 6178
rect 9354 6025 9364 6178
rect 9430 6025 9440 6178
rect 9546 6025 9556 6178
rect 9622 6025 9632 6178
rect 9738 6025 9748 6178
rect 9814 6025 9824 6178
rect 9930 6025 9940 6178
rect 10006 6025 10016 6178
rect 10122 6025 10132 6178
rect 10198 6025 10208 6178
rect 10314 6025 10324 6178
rect 10390 6025 10400 6178
rect 10506 6025 10516 6178
rect 10582 6025 10592 6178
rect 10628 5965 10848 6212
rect 10990 6025 11000 6178
rect 11066 6025 11076 6178
rect 11182 6025 11192 6178
rect 11258 6025 11268 6178
rect 11374 6025 11384 6178
rect 11450 6025 11460 6178
rect 11566 6025 11576 6178
rect 11642 6025 11652 6178
rect 11758 6025 11768 6178
rect 11834 6025 11844 6178
rect 11950 6025 11960 6178
rect 12026 6025 12036 6178
rect 12142 6025 12152 6178
rect 12218 6025 12228 6178
rect 12334 6025 12344 6178
rect 12410 6025 12420 6178
rect 12456 5965 12676 6212
rect 12818 6025 12828 6178
rect 12894 6025 12904 6178
rect 13010 6025 13020 6178
rect 13086 6025 13096 6178
rect 13202 6025 13212 6178
rect 13278 6025 13288 6178
rect 13394 6025 13404 6178
rect 13470 6025 13480 6178
rect 13586 6025 13596 6178
rect 13662 6025 13672 6178
rect 13778 6025 13788 6178
rect 13854 6025 13864 6178
rect 13970 6025 13980 6178
rect 14046 6025 14056 6178
rect 14162 6025 14172 6178
rect 14238 6025 14248 6178
rect 14284 5965 14504 6212
rect 14646 6025 14656 6178
rect 14722 6025 14732 6178
rect 14838 6025 14848 6178
rect 14914 6025 14924 6178
rect 15030 6025 15040 6178
rect 15106 6025 15116 6178
rect 15222 6025 15232 6178
rect 15298 6025 15308 6178
rect 15414 6025 15424 6178
rect 15490 6025 15500 6178
rect 15606 6025 15616 6178
rect 15682 6025 15692 6178
rect 15798 6025 15808 6178
rect 15874 6025 15884 6178
rect 15990 6025 16000 6178
rect 16066 6025 16076 6178
rect 16112 5965 16332 6212
rect 16474 6025 16484 6178
rect 16550 6025 16560 6178
rect 16666 6025 16676 6178
rect 16742 6025 16752 6178
rect 16858 6025 16868 6178
rect 16934 6025 16944 6178
rect 17050 6025 17060 6178
rect 17126 6025 17136 6178
rect 17242 6025 17252 6178
rect 17318 6025 17328 6178
rect 17434 6025 17444 6178
rect 17510 6025 17520 6178
rect 17626 6025 17636 6178
rect 17702 6025 17712 6178
rect 17818 6025 17828 6178
rect 17894 6025 17904 6178
rect 17940 5965 18160 6212
rect 18302 6025 18312 6178
rect 18378 6025 18388 6178
rect 18494 6025 18504 6178
rect 18570 6025 18580 6178
rect 18686 6025 18696 6178
rect 18762 6025 18772 6178
rect 18878 6025 18888 6178
rect 18954 6025 18964 6178
rect 19070 6025 19080 6178
rect 19146 6025 19156 6178
rect 19262 6025 19272 6178
rect 19338 6025 19348 6178
rect 19454 6025 19464 6178
rect 19530 6025 19540 6178
rect 19646 6025 19656 6178
rect 19722 6025 19732 6178
rect 19768 5965 19988 6212
rect 20130 6025 20140 6178
rect 20206 6025 20216 6178
rect 20322 6025 20332 6178
rect 20398 6025 20408 6178
rect 20514 6025 20524 6178
rect 20590 6025 20600 6178
rect 20706 6025 20716 6178
rect 20782 6025 20792 6178
rect 20898 6025 20908 6178
rect 20974 6025 20984 6178
rect 21090 6025 21100 6178
rect 21166 6025 21176 6178
rect 21282 6025 21292 6178
rect 21358 6025 21368 6178
rect 21474 6025 21484 6178
rect 21550 6025 21560 6178
rect 21596 5965 21816 6212
rect 118 5812 128 5965
rect 194 5812 204 5965
rect 310 5812 320 5965
rect 386 5812 396 5965
rect 502 5812 512 5965
rect 578 5812 588 5965
rect 694 5812 704 5965
rect 770 5812 780 5965
rect 886 5812 896 5965
rect 962 5812 972 5965
rect 1078 5812 1088 5965
rect 1154 5812 1164 5965
rect 1270 5812 1280 5965
rect 1346 5812 1356 5965
rect 1462 5812 1472 5965
rect 1528 5812 1708 5965
rect 1946 5812 1956 5965
rect 2022 5812 2032 5965
rect 2138 5812 2148 5965
rect 2214 5812 2224 5965
rect 2330 5812 2340 5965
rect 2406 5812 2416 5965
rect 2522 5812 2532 5965
rect 2598 5812 2608 5965
rect 2714 5812 2724 5965
rect 2790 5812 2800 5965
rect 2906 5812 2916 5965
rect 2982 5812 2992 5965
rect 3098 5812 3108 5965
rect 3174 5812 3184 5965
rect 3290 5812 3300 5965
rect 3356 5812 3536 5965
rect 3774 5812 3784 5965
rect 3850 5812 3860 5965
rect 3966 5812 3976 5965
rect 4042 5812 4052 5965
rect 4158 5812 4168 5965
rect 4234 5812 4244 5965
rect 4350 5812 4360 5965
rect 4426 5812 4436 5965
rect 4542 5812 4552 5965
rect 4618 5812 4628 5965
rect 4734 5812 4744 5965
rect 4810 5812 4820 5965
rect 4926 5812 4936 5965
rect 5002 5812 5012 5965
rect 5118 5812 5128 5965
rect 5184 5812 5364 5965
rect 5602 5812 5612 5965
rect 5678 5812 5688 5965
rect 5794 5812 5804 5965
rect 5870 5812 5880 5965
rect 5986 5812 5996 5965
rect 6062 5812 6072 5965
rect 6178 5812 6188 5965
rect 6254 5812 6264 5965
rect 6370 5812 6380 5965
rect 6446 5812 6456 5965
rect 6562 5812 6572 5965
rect 6638 5812 6648 5965
rect 6754 5812 6764 5965
rect 6830 5812 6840 5965
rect 6946 5812 6956 5965
rect 7012 5812 7192 5965
rect 7430 5812 7440 5965
rect 7506 5812 7516 5965
rect 7622 5812 7632 5965
rect 7698 5812 7708 5965
rect 7814 5812 7824 5965
rect 7890 5812 7900 5965
rect 8006 5812 8016 5965
rect 8082 5812 8092 5965
rect 8198 5812 8208 5965
rect 8274 5812 8284 5965
rect 8390 5812 8400 5965
rect 8466 5812 8476 5965
rect 8582 5812 8592 5965
rect 8658 5812 8668 5965
rect 8774 5812 8784 5965
rect 8840 5812 9020 5965
rect 9258 5812 9268 5965
rect 9334 5812 9344 5965
rect 9450 5812 9460 5965
rect 9526 5812 9536 5965
rect 9642 5812 9652 5965
rect 9718 5812 9728 5965
rect 9834 5812 9844 5965
rect 9910 5812 9920 5965
rect 10026 5812 10036 5965
rect 10102 5812 10112 5965
rect 10218 5812 10228 5965
rect 10294 5812 10304 5965
rect 10410 5812 10420 5965
rect 10486 5812 10496 5965
rect 10602 5812 10612 5965
rect 10668 5812 10848 5965
rect 11086 5812 11096 5965
rect 11162 5812 11172 5965
rect 11278 5812 11288 5965
rect 11354 5812 11364 5965
rect 11470 5812 11480 5965
rect 11546 5812 11556 5965
rect 11662 5812 11672 5965
rect 11738 5812 11748 5965
rect 11854 5812 11864 5965
rect 11930 5812 11940 5965
rect 12046 5812 12056 5965
rect 12122 5812 12132 5965
rect 12238 5812 12248 5965
rect 12314 5812 12324 5965
rect 12430 5812 12440 5965
rect 12496 5812 12676 5965
rect 12914 5812 12924 5965
rect 12990 5812 13000 5965
rect 13106 5812 13116 5965
rect 13182 5812 13192 5965
rect 13298 5812 13308 5965
rect 13374 5812 13384 5965
rect 13490 5812 13500 5965
rect 13566 5812 13576 5965
rect 13682 5812 13692 5965
rect 13758 5812 13768 5965
rect 13874 5812 13884 5965
rect 13950 5812 13960 5965
rect 14066 5812 14076 5965
rect 14142 5812 14152 5965
rect 14258 5812 14268 5965
rect 14324 5812 14504 5965
rect 14742 5812 14752 5965
rect 14818 5812 14828 5965
rect 14934 5812 14944 5965
rect 15010 5812 15020 5965
rect 15126 5812 15136 5965
rect 15202 5812 15212 5965
rect 15318 5812 15328 5965
rect 15394 5812 15404 5965
rect 15510 5812 15520 5965
rect 15586 5812 15596 5965
rect 15702 5812 15712 5965
rect 15778 5812 15788 5965
rect 15894 5812 15904 5965
rect 15970 5812 15980 5965
rect 16086 5812 16096 5965
rect 16152 5812 16332 5965
rect 16570 5812 16580 5965
rect 16646 5812 16656 5965
rect 16762 5812 16772 5965
rect 16838 5812 16848 5965
rect 16954 5812 16964 5965
rect 17030 5812 17040 5965
rect 17146 5812 17156 5965
rect 17222 5812 17232 5965
rect 17338 5812 17348 5965
rect 17414 5812 17424 5965
rect 17530 5812 17540 5965
rect 17606 5812 17616 5965
rect 17722 5812 17732 5965
rect 17798 5812 17808 5965
rect 17914 5812 17924 5965
rect 17980 5812 18160 5965
rect 18398 5812 18408 5965
rect 18474 5812 18484 5965
rect 18590 5812 18600 5965
rect 18666 5812 18676 5965
rect 18782 5812 18792 5965
rect 18858 5812 18868 5965
rect 18974 5812 18984 5965
rect 19050 5812 19060 5965
rect 19166 5812 19176 5965
rect 19242 5812 19252 5965
rect 19358 5812 19368 5965
rect 19434 5812 19444 5965
rect 19550 5812 19560 5965
rect 19626 5812 19636 5965
rect 19742 5812 19752 5965
rect 19808 5812 19988 5965
rect 20226 5812 20236 5965
rect 20302 5812 20312 5965
rect 20418 5812 20428 5965
rect 20494 5812 20504 5965
rect 20610 5812 20620 5965
rect 20686 5812 20696 5965
rect 20802 5812 20812 5965
rect 20878 5812 20888 5965
rect 20994 5812 21004 5965
rect 21070 5812 21080 5965
rect 21186 5812 21196 5965
rect 21262 5812 21272 5965
rect 21378 5812 21388 5965
rect 21454 5812 21464 5965
rect 21570 5812 21580 5965
rect 21636 5812 21816 5965
rect 0 5715 1490 5774
rect 1828 5715 3318 5774
rect 3656 5715 5146 5774
rect 5484 5715 6974 5774
rect 7312 5715 8802 5774
rect 9140 5715 10630 5774
rect 10968 5715 12458 5774
rect 12796 5715 14286 5774
rect 14624 5715 16114 5774
rect 16452 5715 17942 5774
rect 18280 5715 19770 5774
rect 20108 5715 21598 5774
rect 0 5536 1490 5595
rect 1828 5536 3318 5595
rect 3656 5536 5146 5595
rect 5484 5536 6974 5595
rect 7312 5536 8802 5595
rect 9140 5536 10630 5595
rect 10968 5536 12458 5595
rect 12796 5536 14286 5595
rect 14624 5536 16114 5595
rect 16452 5536 17942 5595
rect 18280 5536 19770 5595
rect 20108 5536 21598 5595
rect 22 5311 32 5464
rect 98 5311 108 5464
rect 214 5311 224 5464
rect 290 5311 300 5464
rect 406 5311 416 5464
rect 482 5311 492 5464
rect 598 5311 608 5464
rect 674 5311 684 5464
rect 790 5311 800 5464
rect 866 5311 876 5464
rect 982 5311 992 5464
rect 1058 5311 1068 5464
rect 1174 5311 1184 5464
rect 1250 5311 1260 5464
rect 1366 5311 1376 5464
rect 1442 5311 1452 5464
rect 1488 5251 1708 5498
rect 1850 5311 1860 5464
rect 1926 5311 1936 5464
rect 2042 5311 2052 5464
rect 2118 5311 2128 5464
rect 2234 5311 2244 5464
rect 2310 5311 2320 5464
rect 2426 5311 2436 5464
rect 2502 5311 2512 5464
rect 2618 5311 2628 5464
rect 2694 5311 2704 5464
rect 2810 5311 2820 5464
rect 2886 5311 2896 5464
rect 3002 5311 3012 5464
rect 3078 5311 3088 5464
rect 3194 5311 3204 5464
rect 3270 5311 3280 5464
rect 3316 5251 3536 5498
rect 3678 5311 3688 5464
rect 3754 5311 3764 5464
rect 3870 5311 3880 5464
rect 3946 5311 3956 5464
rect 4062 5311 4072 5464
rect 4138 5311 4148 5464
rect 4254 5311 4264 5464
rect 4330 5311 4340 5464
rect 4446 5311 4456 5464
rect 4522 5311 4532 5464
rect 4638 5311 4648 5464
rect 4714 5311 4724 5464
rect 4830 5311 4840 5464
rect 4906 5311 4916 5464
rect 5022 5311 5032 5464
rect 5098 5311 5108 5464
rect 5144 5251 5364 5498
rect 5506 5311 5516 5464
rect 5582 5311 5592 5464
rect 5698 5311 5708 5464
rect 5774 5311 5784 5464
rect 5890 5311 5900 5464
rect 5966 5311 5976 5464
rect 6082 5311 6092 5464
rect 6158 5311 6168 5464
rect 6274 5311 6284 5464
rect 6350 5311 6360 5464
rect 6466 5311 6476 5464
rect 6542 5311 6552 5464
rect 6658 5311 6668 5464
rect 6734 5311 6744 5464
rect 6850 5311 6860 5464
rect 6926 5311 6936 5464
rect 6972 5251 7192 5498
rect 7334 5311 7344 5464
rect 7410 5311 7420 5464
rect 7526 5311 7536 5464
rect 7602 5311 7612 5464
rect 7718 5311 7728 5464
rect 7794 5311 7804 5464
rect 7910 5311 7920 5464
rect 7986 5311 7996 5464
rect 8102 5311 8112 5464
rect 8178 5311 8188 5464
rect 8294 5311 8304 5464
rect 8370 5311 8380 5464
rect 8486 5311 8496 5464
rect 8562 5311 8572 5464
rect 8678 5311 8688 5464
rect 8754 5311 8764 5464
rect 8800 5251 9020 5498
rect 9162 5311 9172 5464
rect 9238 5311 9248 5464
rect 9354 5311 9364 5464
rect 9430 5311 9440 5464
rect 9546 5311 9556 5464
rect 9622 5311 9632 5464
rect 9738 5311 9748 5464
rect 9814 5311 9824 5464
rect 9930 5311 9940 5464
rect 10006 5311 10016 5464
rect 10122 5311 10132 5464
rect 10198 5311 10208 5464
rect 10314 5311 10324 5464
rect 10390 5311 10400 5464
rect 10506 5311 10516 5464
rect 10582 5311 10592 5464
rect 10628 5251 10848 5498
rect 10990 5311 11000 5464
rect 11066 5311 11076 5464
rect 11182 5311 11192 5464
rect 11258 5311 11268 5464
rect 11374 5311 11384 5464
rect 11450 5311 11460 5464
rect 11566 5311 11576 5464
rect 11642 5311 11652 5464
rect 11758 5311 11768 5464
rect 11834 5311 11844 5464
rect 11950 5311 11960 5464
rect 12026 5311 12036 5464
rect 12142 5311 12152 5464
rect 12218 5311 12228 5464
rect 12334 5311 12344 5464
rect 12410 5311 12420 5464
rect 12456 5251 12676 5498
rect 12818 5311 12828 5464
rect 12894 5311 12904 5464
rect 13010 5311 13020 5464
rect 13086 5311 13096 5464
rect 13202 5311 13212 5464
rect 13278 5311 13288 5464
rect 13394 5311 13404 5464
rect 13470 5311 13480 5464
rect 13586 5311 13596 5464
rect 13662 5311 13672 5464
rect 13778 5311 13788 5464
rect 13854 5311 13864 5464
rect 13970 5311 13980 5464
rect 14046 5311 14056 5464
rect 14162 5311 14172 5464
rect 14238 5311 14248 5464
rect 14284 5251 14504 5498
rect 14646 5311 14656 5464
rect 14722 5311 14732 5464
rect 14838 5311 14848 5464
rect 14914 5311 14924 5464
rect 15030 5311 15040 5464
rect 15106 5311 15116 5464
rect 15222 5311 15232 5464
rect 15298 5311 15308 5464
rect 15414 5311 15424 5464
rect 15490 5311 15500 5464
rect 15606 5311 15616 5464
rect 15682 5311 15692 5464
rect 15798 5311 15808 5464
rect 15874 5311 15884 5464
rect 15990 5311 16000 5464
rect 16066 5311 16076 5464
rect 16112 5251 16332 5498
rect 16474 5311 16484 5464
rect 16550 5311 16560 5464
rect 16666 5311 16676 5464
rect 16742 5311 16752 5464
rect 16858 5311 16868 5464
rect 16934 5311 16944 5464
rect 17050 5311 17060 5464
rect 17126 5311 17136 5464
rect 17242 5311 17252 5464
rect 17318 5311 17328 5464
rect 17434 5311 17444 5464
rect 17510 5311 17520 5464
rect 17626 5311 17636 5464
rect 17702 5311 17712 5464
rect 17818 5311 17828 5464
rect 17894 5311 17904 5464
rect 17940 5251 18160 5498
rect 18302 5311 18312 5464
rect 18378 5311 18388 5464
rect 18494 5311 18504 5464
rect 18570 5311 18580 5464
rect 18686 5311 18696 5464
rect 18762 5311 18772 5464
rect 18878 5311 18888 5464
rect 18954 5311 18964 5464
rect 19070 5311 19080 5464
rect 19146 5311 19156 5464
rect 19262 5311 19272 5464
rect 19338 5311 19348 5464
rect 19454 5311 19464 5464
rect 19530 5311 19540 5464
rect 19646 5311 19656 5464
rect 19722 5311 19732 5464
rect 19768 5251 19988 5498
rect 20130 5311 20140 5464
rect 20206 5311 20216 5464
rect 20322 5311 20332 5464
rect 20398 5311 20408 5464
rect 20514 5311 20524 5464
rect 20590 5311 20600 5464
rect 20706 5311 20716 5464
rect 20782 5311 20792 5464
rect 20898 5311 20908 5464
rect 20974 5311 20984 5464
rect 21090 5311 21100 5464
rect 21166 5311 21176 5464
rect 21282 5311 21292 5464
rect 21358 5311 21368 5464
rect 21474 5311 21484 5464
rect 21550 5311 21560 5464
rect 21596 5251 21816 5498
rect 118 5098 128 5251
rect 194 5098 204 5251
rect 310 5098 320 5251
rect 386 5098 396 5251
rect 502 5098 512 5251
rect 578 5098 588 5251
rect 694 5098 704 5251
rect 770 5098 780 5251
rect 886 5098 896 5251
rect 962 5098 972 5251
rect 1078 5098 1088 5251
rect 1154 5098 1164 5251
rect 1270 5098 1280 5251
rect 1346 5098 1356 5251
rect 1462 5098 1472 5251
rect 1528 5098 1708 5251
rect 1946 5098 1956 5251
rect 2022 5098 2032 5251
rect 2138 5098 2148 5251
rect 2214 5098 2224 5251
rect 2330 5098 2340 5251
rect 2406 5098 2416 5251
rect 2522 5098 2532 5251
rect 2598 5098 2608 5251
rect 2714 5098 2724 5251
rect 2790 5098 2800 5251
rect 2906 5098 2916 5251
rect 2982 5098 2992 5251
rect 3098 5098 3108 5251
rect 3174 5098 3184 5251
rect 3290 5098 3300 5251
rect 3356 5098 3536 5251
rect 3774 5098 3784 5251
rect 3850 5098 3860 5251
rect 3966 5098 3976 5251
rect 4042 5098 4052 5251
rect 4158 5098 4168 5251
rect 4234 5098 4244 5251
rect 4350 5098 4360 5251
rect 4426 5098 4436 5251
rect 4542 5098 4552 5251
rect 4618 5098 4628 5251
rect 4734 5098 4744 5251
rect 4810 5098 4820 5251
rect 4926 5098 4936 5251
rect 5002 5098 5012 5251
rect 5118 5098 5128 5251
rect 5184 5098 5364 5251
rect 5602 5098 5612 5251
rect 5678 5098 5688 5251
rect 5794 5098 5804 5251
rect 5870 5098 5880 5251
rect 5986 5098 5996 5251
rect 6062 5098 6072 5251
rect 6178 5098 6188 5251
rect 6254 5098 6264 5251
rect 6370 5098 6380 5251
rect 6446 5098 6456 5251
rect 6562 5098 6572 5251
rect 6638 5098 6648 5251
rect 6754 5098 6764 5251
rect 6830 5098 6840 5251
rect 6946 5098 6956 5251
rect 7012 5098 7192 5251
rect 7430 5098 7440 5251
rect 7506 5098 7516 5251
rect 7622 5098 7632 5251
rect 7698 5098 7708 5251
rect 7814 5098 7824 5251
rect 7890 5098 7900 5251
rect 8006 5098 8016 5251
rect 8082 5098 8092 5251
rect 8198 5098 8208 5251
rect 8274 5098 8284 5251
rect 8390 5098 8400 5251
rect 8466 5098 8476 5251
rect 8582 5098 8592 5251
rect 8658 5098 8668 5251
rect 8774 5098 8784 5251
rect 8840 5098 9020 5251
rect 9258 5098 9268 5251
rect 9334 5098 9344 5251
rect 9450 5098 9460 5251
rect 9526 5098 9536 5251
rect 9642 5098 9652 5251
rect 9718 5098 9728 5251
rect 9834 5098 9844 5251
rect 9910 5098 9920 5251
rect 10026 5098 10036 5251
rect 10102 5098 10112 5251
rect 10218 5098 10228 5251
rect 10294 5098 10304 5251
rect 10410 5098 10420 5251
rect 10486 5098 10496 5251
rect 10602 5098 10612 5251
rect 10668 5098 10848 5251
rect 11086 5098 11096 5251
rect 11162 5098 11172 5251
rect 11278 5098 11288 5251
rect 11354 5098 11364 5251
rect 11470 5098 11480 5251
rect 11546 5098 11556 5251
rect 11662 5098 11672 5251
rect 11738 5098 11748 5251
rect 11854 5098 11864 5251
rect 11930 5098 11940 5251
rect 12046 5098 12056 5251
rect 12122 5098 12132 5251
rect 12238 5098 12248 5251
rect 12314 5098 12324 5251
rect 12430 5098 12440 5251
rect 12496 5098 12676 5251
rect 12914 5098 12924 5251
rect 12990 5098 13000 5251
rect 13106 5098 13116 5251
rect 13182 5098 13192 5251
rect 13298 5098 13308 5251
rect 13374 5098 13384 5251
rect 13490 5098 13500 5251
rect 13566 5098 13576 5251
rect 13682 5098 13692 5251
rect 13758 5098 13768 5251
rect 13874 5098 13884 5251
rect 13950 5098 13960 5251
rect 14066 5098 14076 5251
rect 14142 5098 14152 5251
rect 14258 5098 14268 5251
rect 14324 5098 14504 5251
rect 14742 5098 14752 5251
rect 14818 5098 14828 5251
rect 14934 5098 14944 5251
rect 15010 5098 15020 5251
rect 15126 5098 15136 5251
rect 15202 5098 15212 5251
rect 15318 5098 15328 5251
rect 15394 5098 15404 5251
rect 15510 5098 15520 5251
rect 15586 5098 15596 5251
rect 15702 5098 15712 5251
rect 15778 5098 15788 5251
rect 15894 5098 15904 5251
rect 15970 5098 15980 5251
rect 16086 5098 16096 5251
rect 16152 5098 16332 5251
rect 16570 5098 16580 5251
rect 16646 5098 16656 5251
rect 16762 5098 16772 5251
rect 16838 5098 16848 5251
rect 16954 5098 16964 5251
rect 17030 5098 17040 5251
rect 17146 5098 17156 5251
rect 17222 5098 17232 5251
rect 17338 5098 17348 5251
rect 17414 5098 17424 5251
rect 17530 5098 17540 5251
rect 17606 5098 17616 5251
rect 17722 5098 17732 5251
rect 17798 5098 17808 5251
rect 17914 5098 17924 5251
rect 17980 5098 18160 5251
rect 18398 5098 18408 5251
rect 18474 5098 18484 5251
rect 18590 5098 18600 5251
rect 18666 5098 18676 5251
rect 18782 5098 18792 5251
rect 18858 5098 18868 5251
rect 18974 5098 18984 5251
rect 19050 5098 19060 5251
rect 19166 5098 19176 5251
rect 19242 5098 19252 5251
rect 19358 5098 19368 5251
rect 19434 5098 19444 5251
rect 19550 5098 19560 5251
rect 19626 5098 19636 5251
rect 19742 5098 19752 5251
rect 19808 5098 19988 5251
rect 20226 5098 20236 5251
rect 20302 5098 20312 5251
rect 20418 5098 20428 5251
rect 20494 5098 20504 5251
rect 20610 5098 20620 5251
rect 20686 5098 20696 5251
rect 20802 5098 20812 5251
rect 20878 5098 20888 5251
rect 20994 5098 21004 5251
rect 21070 5098 21080 5251
rect 21186 5098 21196 5251
rect 21262 5098 21272 5251
rect 21378 5098 21388 5251
rect 21454 5098 21464 5251
rect 21570 5098 21580 5251
rect 21636 5098 21816 5251
rect 0 5001 1490 5060
rect 1828 5001 3318 5060
rect 3656 5001 5146 5060
rect 5484 5001 6974 5060
rect 7312 5001 8802 5060
rect 9140 5001 10630 5060
rect 10968 5001 12458 5060
rect 12796 5001 14286 5060
rect 14624 5001 16114 5060
rect 16452 5001 17942 5060
rect 18280 5001 19770 5060
rect 20108 5001 21598 5060
rect 0 4822 1490 4881
rect 1828 4822 3318 4881
rect 3656 4822 5146 4881
rect 5484 4822 6974 4881
rect 7312 4822 8802 4881
rect 9140 4822 10630 4881
rect 10968 4822 12458 4881
rect 12796 4822 14286 4881
rect 14624 4822 16114 4881
rect 16452 4822 17942 4881
rect 18280 4822 19770 4881
rect 20108 4822 21598 4881
rect 22 4597 32 4750
rect 98 4597 108 4750
rect 214 4597 224 4750
rect 290 4597 300 4750
rect 406 4597 416 4750
rect 482 4597 492 4750
rect 598 4597 608 4750
rect 674 4597 684 4750
rect 790 4597 800 4750
rect 866 4597 876 4750
rect 982 4597 992 4750
rect 1058 4597 1068 4750
rect 1174 4597 1184 4750
rect 1250 4597 1260 4750
rect 1366 4597 1376 4750
rect 1442 4597 1452 4750
rect 1488 4537 1708 4784
rect 1850 4597 1860 4750
rect 1926 4597 1936 4750
rect 2042 4597 2052 4750
rect 2118 4597 2128 4750
rect 2234 4597 2244 4750
rect 2310 4597 2320 4750
rect 2426 4597 2436 4750
rect 2502 4597 2512 4750
rect 2618 4597 2628 4750
rect 2694 4597 2704 4750
rect 2810 4597 2820 4750
rect 2886 4597 2896 4750
rect 3002 4597 3012 4750
rect 3078 4597 3088 4750
rect 3194 4597 3204 4750
rect 3270 4597 3280 4750
rect 3316 4537 3536 4784
rect 3678 4597 3688 4750
rect 3754 4597 3764 4750
rect 3870 4597 3880 4750
rect 3946 4597 3956 4750
rect 4062 4597 4072 4750
rect 4138 4597 4148 4750
rect 4254 4597 4264 4750
rect 4330 4597 4340 4750
rect 4446 4597 4456 4750
rect 4522 4597 4532 4750
rect 4638 4597 4648 4750
rect 4714 4597 4724 4750
rect 4830 4597 4840 4750
rect 4906 4597 4916 4750
rect 5022 4597 5032 4750
rect 5098 4597 5108 4750
rect 5144 4537 5364 4784
rect 5506 4597 5516 4750
rect 5582 4597 5592 4750
rect 5698 4597 5708 4750
rect 5774 4597 5784 4750
rect 5890 4597 5900 4750
rect 5966 4597 5976 4750
rect 6082 4597 6092 4750
rect 6158 4597 6168 4750
rect 6274 4597 6284 4750
rect 6350 4597 6360 4750
rect 6466 4597 6476 4750
rect 6542 4597 6552 4750
rect 6658 4597 6668 4750
rect 6734 4597 6744 4750
rect 6850 4597 6860 4750
rect 6926 4597 6936 4750
rect 6972 4537 7192 4784
rect 7334 4597 7344 4750
rect 7410 4597 7420 4750
rect 7526 4597 7536 4750
rect 7602 4597 7612 4750
rect 7718 4597 7728 4750
rect 7794 4597 7804 4750
rect 7910 4597 7920 4750
rect 7986 4597 7996 4750
rect 8102 4597 8112 4750
rect 8178 4597 8188 4750
rect 8294 4597 8304 4750
rect 8370 4597 8380 4750
rect 8486 4597 8496 4750
rect 8562 4597 8572 4750
rect 8678 4597 8688 4750
rect 8754 4597 8764 4750
rect 8800 4537 9020 4784
rect 9162 4597 9172 4750
rect 9238 4597 9248 4750
rect 9354 4597 9364 4750
rect 9430 4597 9440 4750
rect 9546 4597 9556 4750
rect 9622 4597 9632 4750
rect 9738 4597 9748 4750
rect 9814 4597 9824 4750
rect 9930 4597 9940 4750
rect 10006 4597 10016 4750
rect 10122 4597 10132 4750
rect 10198 4597 10208 4750
rect 10314 4597 10324 4750
rect 10390 4597 10400 4750
rect 10506 4597 10516 4750
rect 10582 4597 10592 4750
rect 10628 4537 10848 4784
rect 10990 4597 11000 4750
rect 11066 4597 11076 4750
rect 11182 4597 11192 4750
rect 11258 4597 11268 4750
rect 11374 4597 11384 4750
rect 11450 4597 11460 4750
rect 11566 4597 11576 4750
rect 11642 4597 11652 4750
rect 11758 4597 11768 4750
rect 11834 4597 11844 4750
rect 11950 4597 11960 4750
rect 12026 4597 12036 4750
rect 12142 4597 12152 4750
rect 12218 4597 12228 4750
rect 12334 4597 12344 4750
rect 12410 4597 12420 4750
rect 12456 4537 12676 4784
rect 12818 4597 12828 4750
rect 12894 4597 12904 4750
rect 13010 4597 13020 4750
rect 13086 4597 13096 4750
rect 13202 4597 13212 4750
rect 13278 4597 13288 4750
rect 13394 4597 13404 4750
rect 13470 4597 13480 4750
rect 13586 4597 13596 4750
rect 13662 4597 13672 4750
rect 13778 4597 13788 4750
rect 13854 4597 13864 4750
rect 13970 4597 13980 4750
rect 14046 4597 14056 4750
rect 14162 4597 14172 4750
rect 14238 4597 14248 4750
rect 14284 4537 14504 4784
rect 14646 4597 14656 4750
rect 14722 4597 14732 4750
rect 14838 4597 14848 4750
rect 14914 4597 14924 4750
rect 15030 4597 15040 4750
rect 15106 4597 15116 4750
rect 15222 4597 15232 4750
rect 15298 4597 15308 4750
rect 15414 4597 15424 4750
rect 15490 4597 15500 4750
rect 15606 4597 15616 4750
rect 15682 4597 15692 4750
rect 15798 4597 15808 4750
rect 15874 4597 15884 4750
rect 15990 4597 16000 4750
rect 16066 4597 16076 4750
rect 16112 4537 16332 4784
rect 16474 4597 16484 4750
rect 16550 4597 16560 4750
rect 16666 4597 16676 4750
rect 16742 4597 16752 4750
rect 16858 4597 16868 4750
rect 16934 4597 16944 4750
rect 17050 4597 17060 4750
rect 17126 4597 17136 4750
rect 17242 4597 17252 4750
rect 17318 4597 17328 4750
rect 17434 4597 17444 4750
rect 17510 4597 17520 4750
rect 17626 4597 17636 4750
rect 17702 4597 17712 4750
rect 17818 4597 17828 4750
rect 17894 4597 17904 4750
rect 17940 4537 18160 4784
rect 18302 4597 18312 4750
rect 18378 4597 18388 4750
rect 18494 4597 18504 4750
rect 18570 4597 18580 4750
rect 18686 4597 18696 4750
rect 18762 4597 18772 4750
rect 18878 4597 18888 4750
rect 18954 4597 18964 4750
rect 19070 4597 19080 4750
rect 19146 4597 19156 4750
rect 19262 4597 19272 4750
rect 19338 4597 19348 4750
rect 19454 4597 19464 4750
rect 19530 4597 19540 4750
rect 19646 4597 19656 4750
rect 19722 4597 19732 4750
rect 19768 4537 19988 4784
rect 20130 4597 20140 4750
rect 20206 4597 20216 4750
rect 20322 4597 20332 4750
rect 20398 4597 20408 4750
rect 20514 4597 20524 4750
rect 20590 4597 20600 4750
rect 20706 4597 20716 4750
rect 20782 4597 20792 4750
rect 20898 4597 20908 4750
rect 20974 4597 20984 4750
rect 21090 4597 21100 4750
rect 21166 4597 21176 4750
rect 21282 4597 21292 4750
rect 21358 4597 21368 4750
rect 21474 4597 21484 4750
rect 21550 4597 21560 4750
rect 21596 4537 21816 4784
rect 118 4384 128 4537
rect 194 4384 204 4537
rect 310 4384 320 4537
rect 386 4384 396 4537
rect 502 4384 512 4537
rect 578 4384 588 4537
rect 694 4384 704 4537
rect 770 4384 780 4537
rect 886 4384 896 4537
rect 962 4384 972 4537
rect 1078 4384 1088 4537
rect 1154 4384 1164 4537
rect 1270 4384 1280 4537
rect 1346 4384 1356 4537
rect 1462 4384 1472 4537
rect 1528 4384 1708 4537
rect 1946 4384 1956 4537
rect 2022 4384 2032 4537
rect 2138 4384 2148 4537
rect 2214 4384 2224 4537
rect 2330 4384 2340 4537
rect 2406 4384 2416 4537
rect 2522 4384 2532 4537
rect 2598 4384 2608 4537
rect 2714 4384 2724 4537
rect 2790 4384 2800 4537
rect 2906 4384 2916 4537
rect 2982 4384 2992 4537
rect 3098 4384 3108 4537
rect 3174 4384 3184 4537
rect 3290 4384 3300 4537
rect 3356 4384 3536 4537
rect 3774 4384 3784 4537
rect 3850 4384 3860 4537
rect 3966 4384 3976 4537
rect 4042 4384 4052 4537
rect 4158 4384 4168 4537
rect 4234 4384 4244 4537
rect 4350 4384 4360 4537
rect 4426 4384 4436 4537
rect 4542 4384 4552 4537
rect 4618 4384 4628 4537
rect 4734 4384 4744 4537
rect 4810 4384 4820 4537
rect 4926 4384 4936 4537
rect 5002 4384 5012 4537
rect 5118 4384 5128 4537
rect 5184 4384 5364 4537
rect 5602 4384 5612 4537
rect 5678 4384 5688 4537
rect 5794 4384 5804 4537
rect 5870 4384 5880 4537
rect 5986 4384 5996 4537
rect 6062 4384 6072 4537
rect 6178 4384 6188 4537
rect 6254 4384 6264 4537
rect 6370 4384 6380 4537
rect 6446 4384 6456 4537
rect 6562 4384 6572 4537
rect 6638 4384 6648 4537
rect 6754 4384 6764 4537
rect 6830 4384 6840 4537
rect 6946 4384 6956 4537
rect 7012 4384 7192 4537
rect 7430 4384 7440 4537
rect 7506 4384 7516 4537
rect 7622 4384 7632 4537
rect 7698 4384 7708 4537
rect 7814 4384 7824 4537
rect 7890 4384 7900 4537
rect 8006 4384 8016 4537
rect 8082 4384 8092 4537
rect 8198 4384 8208 4537
rect 8274 4384 8284 4537
rect 8390 4384 8400 4537
rect 8466 4384 8476 4537
rect 8582 4384 8592 4537
rect 8658 4384 8668 4537
rect 8774 4384 8784 4537
rect 8840 4384 9020 4537
rect 9258 4384 9268 4537
rect 9334 4384 9344 4537
rect 9450 4384 9460 4537
rect 9526 4384 9536 4537
rect 9642 4384 9652 4537
rect 9718 4384 9728 4537
rect 9834 4384 9844 4537
rect 9910 4384 9920 4537
rect 10026 4384 10036 4537
rect 10102 4384 10112 4537
rect 10218 4384 10228 4537
rect 10294 4384 10304 4537
rect 10410 4384 10420 4537
rect 10486 4384 10496 4537
rect 10602 4384 10612 4537
rect 10668 4384 10848 4537
rect 11086 4384 11096 4537
rect 11162 4384 11172 4537
rect 11278 4384 11288 4537
rect 11354 4384 11364 4537
rect 11470 4384 11480 4537
rect 11546 4384 11556 4537
rect 11662 4384 11672 4537
rect 11738 4384 11748 4537
rect 11854 4384 11864 4537
rect 11930 4384 11940 4537
rect 12046 4384 12056 4537
rect 12122 4384 12132 4537
rect 12238 4384 12248 4537
rect 12314 4384 12324 4537
rect 12430 4384 12440 4537
rect 12496 4384 12676 4537
rect 12914 4384 12924 4537
rect 12990 4384 13000 4537
rect 13106 4384 13116 4537
rect 13182 4384 13192 4537
rect 13298 4384 13308 4537
rect 13374 4384 13384 4537
rect 13490 4384 13500 4537
rect 13566 4384 13576 4537
rect 13682 4384 13692 4537
rect 13758 4384 13768 4537
rect 13874 4384 13884 4537
rect 13950 4384 13960 4537
rect 14066 4384 14076 4537
rect 14142 4384 14152 4537
rect 14258 4384 14268 4537
rect 14324 4384 14504 4537
rect 14742 4384 14752 4537
rect 14818 4384 14828 4537
rect 14934 4384 14944 4537
rect 15010 4384 15020 4537
rect 15126 4384 15136 4537
rect 15202 4384 15212 4537
rect 15318 4384 15328 4537
rect 15394 4384 15404 4537
rect 15510 4384 15520 4537
rect 15586 4384 15596 4537
rect 15702 4384 15712 4537
rect 15778 4384 15788 4537
rect 15894 4384 15904 4537
rect 15970 4384 15980 4537
rect 16086 4384 16096 4537
rect 16152 4384 16332 4537
rect 16570 4384 16580 4537
rect 16646 4384 16656 4537
rect 16762 4384 16772 4537
rect 16838 4384 16848 4537
rect 16954 4384 16964 4537
rect 17030 4384 17040 4537
rect 17146 4384 17156 4537
rect 17222 4384 17232 4537
rect 17338 4384 17348 4537
rect 17414 4384 17424 4537
rect 17530 4384 17540 4537
rect 17606 4384 17616 4537
rect 17722 4384 17732 4537
rect 17798 4384 17808 4537
rect 17914 4384 17924 4537
rect 17980 4384 18160 4537
rect 18398 4384 18408 4537
rect 18474 4384 18484 4537
rect 18590 4384 18600 4537
rect 18666 4384 18676 4537
rect 18782 4384 18792 4537
rect 18858 4384 18868 4537
rect 18974 4384 18984 4537
rect 19050 4384 19060 4537
rect 19166 4384 19176 4537
rect 19242 4384 19252 4537
rect 19358 4384 19368 4537
rect 19434 4384 19444 4537
rect 19550 4384 19560 4537
rect 19626 4384 19636 4537
rect 19742 4384 19752 4537
rect 19808 4384 19988 4537
rect 20226 4384 20236 4537
rect 20302 4384 20312 4537
rect 20418 4384 20428 4537
rect 20494 4384 20504 4537
rect 20610 4384 20620 4537
rect 20686 4384 20696 4537
rect 20802 4384 20812 4537
rect 20878 4384 20888 4537
rect 20994 4384 21004 4537
rect 21070 4384 21080 4537
rect 21186 4384 21196 4537
rect 21262 4384 21272 4537
rect 21378 4384 21388 4537
rect 21454 4384 21464 4537
rect 21570 4384 21580 4537
rect 21636 4384 21816 4537
rect 0 4287 1490 4346
rect 1828 4287 3318 4346
rect 3656 4287 5146 4346
rect 5484 4287 6974 4346
rect 7312 4287 8802 4346
rect 9140 4287 10630 4346
rect 10968 4287 12458 4346
rect 12796 4287 14286 4346
rect 14624 4287 16114 4346
rect 16452 4287 17942 4346
rect 18280 4287 19770 4346
rect 20108 4287 21598 4346
rect 0 4108 1490 4167
rect 1828 4108 3318 4167
rect 3656 4108 5146 4167
rect 5484 4108 6974 4167
rect 7312 4108 8802 4167
rect 9140 4108 10630 4167
rect 10968 4108 12458 4167
rect 12796 4108 14286 4167
rect 14624 4108 16114 4167
rect 16452 4108 17942 4167
rect 18280 4108 19770 4167
rect 20108 4108 21598 4167
rect 22 3883 32 4036
rect 98 3883 108 4036
rect 214 3883 224 4036
rect 290 3883 300 4036
rect 406 3883 416 4036
rect 482 3883 492 4036
rect 598 3883 608 4036
rect 674 3883 684 4036
rect 790 3883 800 4036
rect 866 3883 876 4036
rect 982 3883 992 4036
rect 1058 3883 1068 4036
rect 1174 3883 1184 4036
rect 1250 3883 1260 4036
rect 1366 3883 1376 4036
rect 1442 3883 1452 4036
rect 1488 3823 1708 4070
rect 1850 3883 1860 4036
rect 1926 3883 1936 4036
rect 2042 3883 2052 4036
rect 2118 3883 2128 4036
rect 2234 3883 2244 4036
rect 2310 3883 2320 4036
rect 2426 3883 2436 4036
rect 2502 3883 2512 4036
rect 2618 3883 2628 4036
rect 2694 3883 2704 4036
rect 2810 3883 2820 4036
rect 2886 3883 2896 4036
rect 3002 3883 3012 4036
rect 3078 3883 3088 4036
rect 3194 3883 3204 4036
rect 3270 3883 3280 4036
rect 3316 3823 3536 4070
rect 3678 3883 3688 4036
rect 3754 3883 3764 4036
rect 3870 3883 3880 4036
rect 3946 3883 3956 4036
rect 4062 3883 4072 4036
rect 4138 3883 4148 4036
rect 4254 3883 4264 4036
rect 4330 3883 4340 4036
rect 4446 3883 4456 4036
rect 4522 3883 4532 4036
rect 4638 3883 4648 4036
rect 4714 3883 4724 4036
rect 4830 3883 4840 4036
rect 4906 3883 4916 4036
rect 5022 3883 5032 4036
rect 5098 3883 5108 4036
rect 5144 3823 5364 4070
rect 5506 3883 5516 4036
rect 5582 3883 5592 4036
rect 5698 3883 5708 4036
rect 5774 3883 5784 4036
rect 5890 3883 5900 4036
rect 5966 3883 5976 4036
rect 6082 3883 6092 4036
rect 6158 3883 6168 4036
rect 6274 3883 6284 4036
rect 6350 3883 6360 4036
rect 6466 3883 6476 4036
rect 6542 3883 6552 4036
rect 6658 3883 6668 4036
rect 6734 3883 6744 4036
rect 6850 3883 6860 4036
rect 6926 3883 6936 4036
rect 6972 3823 7192 4070
rect 7334 3883 7344 4036
rect 7410 3883 7420 4036
rect 7526 3883 7536 4036
rect 7602 3883 7612 4036
rect 7718 3883 7728 4036
rect 7794 3883 7804 4036
rect 7910 3883 7920 4036
rect 7986 3883 7996 4036
rect 8102 3883 8112 4036
rect 8178 3883 8188 4036
rect 8294 3883 8304 4036
rect 8370 3883 8380 4036
rect 8486 3883 8496 4036
rect 8562 3883 8572 4036
rect 8678 3883 8688 4036
rect 8754 3883 8764 4036
rect 8800 3823 9020 4070
rect 9162 3883 9172 4036
rect 9238 3883 9248 4036
rect 9354 3883 9364 4036
rect 9430 3883 9440 4036
rect 9546 3883 9556 4036
rect 9622 3883 9632 4036
rect 9738 3883 9748 4036
rect 9814 3883 9824 4036
rect 9930 3883 9940 4036
rect 10006 3883 10016 4036
rect 10122 3883 10132 4036
rect 10198 3883 10208 4036
rect 10314 3883 10324 4036
rect 10390 3883 10400 4036
rect 10506 3883 10516 4036
rect 10582 3883 10592 4036
rect 10628 3823 10848 4070
rect 10990 3883 11000 4036
rect 11066 3883 11076 4036
rect 11182 3883 11192 4036
rect 11258 3883 11268 4036
rect 11374 3883 11384 4036
rect 11450 3883 11460 4036
rect 11566 3883 11576 4036
rect 11642 3883 11652 4036
rect 11758 3883 11768 4036
rect 11834 3883 11844 4036
rect 11950 3883 11960 4036
rect 12026 3883 12036 4036
rect 12142 3883 12152 4036
rect 12218 3883 12228 4036
rect 12334 3883 12344 4036
rect 12410 3883 12420 4036
rect 12456 3823 12676 4070
rect 12818 3883 12828 4036
rect 12894 3883 12904 4036
rect 13010 3883 13020 4036
rect 13086 3883 13096 4036
rect 13202 3883 13212 4036
rect 13278 3883 13288 4036
rect 13394 3883 13404 4036
rect 13470 3883 13480 4036
rect 13586 3883 13596 4036
rect 13662 3883 13672 4036
rect 13778 3883 13788 4036
rect 13854 3883 13864 4036
rect 13970 3883 13980 4036
rect 14046 3883 14056 4036
rect 14162 3883 14172 4036
rect 14238 3883 14248 4036
rect 14284 3823 14504 4070
rect 14646 3883 14656 4036
rect 14722 3883 14732 4036
rect 14838 3883 14848 4036
rect 14914 3883 14924 4036
rect 15030 3883 15040 4036
rect 15106 3883 15116 4036
rect 15222 3883 15232 4036
rect 15298 3883 15308 4036
rect 15414 3883 15424 4036
rect 15490 3883 15500 4036
rect 15606 3883 15616 4036
rect 15682 3883 15692 4036
rect 15798 3883 15808 4036
rect 15874 3883 15884 4036
rect 15990 3883 16000 4036
rect 16066 3883 16076 4036
rect 16112 3823 16332 4070
rect 16474 3883 16484 4036
rect 16550 3883 16560 4036
rect 16666 3883 16676 4036
rect 16742 3883 16752 4036
rect 16858 3883 16868 4036
rect 16934 3883 16944 4036
rect 17050 3883 17060 4036
rect 17126 3883 17136 4036
rect 17242 3883 17252 4036
rect 17318 3883 17328 4036
rect 17434 3883 17444 4036
rect 17510 3883 17520 4036
rect 17626 3883 17636 4036
rect 17702 3883 17712 4036
rect 17818 3883 17828 4036
rect 17894 3883 17904 4036
rect 17940 3823 18160 4070
rect 18302 3883 18312 4036
rect 18378 3883 18388 4036
rect 18494 3883 18504 4036
rect 18570 3883 18580 4036
rect 18686 3883 18696 4036
rect 18762 3883 18772 4036
rect 18878 3883 18888 4036
rect 18954 3883 18964 4036
rect 19070 3883 19080 4036
rect 19146 3883 19156 4036
rect 19262 3883 19272 4036
rect 19338 3883 19348 4036
rect 19454 3883 19464 4036
rect 19530 3883 19540 4036
rect 19646 3883 19656 4036
rect 19722 3883 19732 4036
rect 19768 3823 19988 4070
rect 20130 3883 20140 4036
rect 20206 3883 20216 4036
rect 20322 3883 20332 4036
rect 20398 3883 20408 4036
rect 20514 3883 20524 4036
rect 20590 3883 20600 4036
rect 20706 3883 20716 4036
rect 20782 3883 20792 4036
rect 20898 3883 20908 4036
rect 20974 3883 20984 4036
rect 21090 3883 21100 4036
rect 21166 3883 21176 4036
rect 21282 3883 21292 4036
rect 21358 3883 21368 4036
rect 21474 3883 21484 4036
rect 21550 3883 21560 4036
rect 21596 3823 21816 4070
rect 118 3670 128 3823
rect 194 3670 204 3823
rect 310 3670 320 3823
rect 386 3670 396 3823
rect 502 3670 512 3823
rect 578 3670 588 3823
rect 694 3670 704 3823
rect 770 3670 780 3823
rect 886 3670 896 3823
rect 962 3670 972 3823
rect 1078 3670 1088 3823
rect 1154 3670 1164 3823
rect 1270 3670 1280 3823
rect 1346 3670 1356 3823
rect 1462 3670 1472 3823
rect 1528 3670 1708 3823
rect 1946 3670 1956 3823
rect 2022 3670 2032 3823
rect 2138 3670 2148 3823
rect 2214 3670 2224 3823
rect 2330 3670 2340 3823
rect 2406 3670 2416 3823
rect 2522 3670 2532 3823
rect 2598 3670 2608 3823
rect 2714 3670 2724 3823
rect 2790 3670 2800 3823
rect 2906 3670 2916 3823
rect 2982 3670 2992 3823
rect 3098 3670 3108 3823
rect 3174 3670 3184 3823
rect 3290 3670 3300 3823
rect 3356 3670 3536 3823
rect 3774 3670 3784 3823
rect 3850 3670 3860 3823
rect 3966 3670 3976 3823
rect 4042 3670 4052 3823
rect 4158 3670 4168 3823
rect 4234 3670 4244 3823
rect 4350 3670 4360 3823
rect 4426 3670 4436 3823
rect 4542 3670 4552 3823
rect 4618 3670 4628 3823
rect 4734 3670 4744 3823
rect 4810 3670 4820 3823
rect 4926 3670 4936 3823
rect 5002 3670 5012 3823
rect 5118 3670 5128 3823
rect 5184 3670 5364 3823
rect 5602 3670 5612 3823
rect 5678 3670 5688 3823
rect 5794 3670 5804 3823
rect 5870 3670 5880 3823
rect 5986 3670 5996 3823
rect 6062 3670 6072 3823
rect 6178 3670 6188 3823
rect 6254 3670 6264 3823
rect 6370 3670 6380 3823
rect 6446 3670 6456 3823
rect 6562 3670 6572 3823
rect 6638 3670 6648 3823
rect 6754 3670 6764 3823
rect 6830 3670 6840 3823
rect 6946 3670 6956 3823
rect 7012 3670 7192 3823
rect 7430 3670 7440 3823
rect 7506 3670 7516 3823
rect 7622 3670 7632 3823
rect 7698 3670 7708 3823
rect 7814 3670 7824 3823
rect 7890 3670 7900 3823
rect 8006 3670 8016 3823
rect 8082 3670 8092 3823
rect 8198 3670 8208 3823
rect 8274 3670 8284 3823
rect 8390 3670 8400 3823
rect 8466 3670 8476 3823
rect 8582 3670 8592 3823
rect 8658 3670 8668 3823
rect 8774 3670 8784 3823
rect 8840 3670 9020 3823
rect 9258 3670 9268 3823
rect 9334 3670 9344 3823
rect 9450 3670 9460 3823
rect 9526 3670 9536 3823
rect 9642 3670 9652 3823
rect 9718 3670 9728 3823
rect 9834 3670 9844 3823
rect 9910 3670 9920 3823
rect 10026 3670 10036 3823
rect 10102 3670 10112 3823
rect 10218 3670 10228 3823
rect 10294 3670 10304 3823
rect 10410 3670 10420 3823
rect 10486 3670 10496 3823
rect 10602 3670 10612 3823
rect 10668 3670 10848 3823
rect 11086 3670 11096 3823
rect 11162 3670 11172 3823
rect 11278 3670 11288 3823
rect 11354 3670 11364 3823
rect 11470 3670 11480 3823
rect 11546 3670 11556 3823
rect 11662 3670 11672 3823
rect 11738 3670 11748 3823
rect 11854 3670 11864 3823
rect 11930 3670 11940 3823
rect 12046 3670 12056 3823
rect 12122 3670 12132 3823
rect 12238 3670 12248 3823
rect 12314 3670 12324 3823
rect 12430 3670 12440 3823
rect 12496 3670 12676 3823
rect 12914 3670 12924 3823
rect 12990 3670 13000 3823
rect 13106 3670 13116 3823
rect 13182 3670 13192 3823
rect 13298 3670 13308 3823
rect 13374 3670 13384 3823
rect 13490 3670 13500 3823
rect 13566 3670 13576 3823
rect 13682 3670 13692 3823
rect 13758 3670 13768 3823
rect 13874 3670 13884 3823
rect 13950 3670 13960 3823
rect 14066 3670 14076 3823
rect 14142 3670 14152 3823
rect 14258 3670 14268 3823
rect 14324 3670 14504 3823
rect 14742 3670 14752 3823
rect 14818 3670 14828 3823
rect 14934 3670 14944 3823
rect 15010 3670 15020 3823
rect 15126 3670 15136 3823
rect 15202 3670 15212 3823
rect 15318 3670 15328 3823
rect 15394 3670 15404 3823
rect 15510 3670 15520 3823
rect 15586 3670 15596 3823
rect 15702 3670 15712 3823
rect 15778 3670 15788 3823
rect 15894 3670 15904 3823
rect 15970 3670 15980 3823
rect 16086 3670 16096 3823
rect 16152 3670 16332 3823
rect 16570 3670 16580 3823
rect 16646 3670 16656 3823
rect 16762 3670 16772 3823
rect 16838 3670 16848 3823
rect 16954 3670 16964 3823
rect 17030 3670 17040 3823
rect 17146 3670 17156 3823
rect 17222 3670 17232 3823
rect 17338 3670 17348 3823
rect 17414 3670 17424 3823
rect 17530 3670 17540 3823
rect 17606 3670 17616 3823
rect 17722 3670 17732 3823
rect 17798 3670 17808 3823
rect 17914 3670 17924 3823
rect 17980 3670 18160 3823
rect 18398 3670 18408 3823
rect 18474 3670 18484 3823
rect 18590 3670 18600 3823
rect 18666 3670 18676 3823
rect 18782 3670 18792 3823
rect 18858 3670 18868 3823
rect 18974 3670 18984 3823
rect 19050 3670 19060 3823
rect 19166 3670 19176 3823
rect 19242 3670 19252 3823
rect 19358 3670 19368 3823
rect 19434 3670 19444 3823
rect 19550 3670 19560 3823
rect 19626 3670 19636 3823
rect 19742 3670 19752 3823
rect 19808 3670 19988 3823
rect 20226 3670 20236 3823
rect 20302 3670 20312 3823
rect 20418 3670 20428 3823
rect 20494 3670 20504 3823
rect 20610 3670 20620 3823
rect 20686 3670 20696 3823
rect 20802 3670 20812 3823
rect 20878 3670 20888 3823
rect 20994 3670 21004 3823
rect 21070 3670 21080 3823
rect 21186 3670 21196 3823
rect 21262 3670 21272 3823
rect 21378 3670 21388 3823
rect 21454 3670 21464 3823
rect 21570 3670 21580 3823
rect 21636 3670 21816 3823
rect 0 3573 1490 3632
rect 1828 3573 3318 3632
rect 3656 3573 5146 3632
rect 5484 3573 6974 3632
rect 7312 3573 8802 3632
rect 9140 3573 10630 3632
rect 10968 3573 12458 3632
rect 12796 3573 14286 3632
rect 14624 3573 16114 3632
rect 16452 3573 17942 3632
rect 18280 3573 19770 3632
rect 20108 3573 21598 3632
rect 0 3394 1490 3453
rect 1828 3394 3318 3453
rect 3656 3394 5146 3453
rect 5484 3394 6974 3453
rect 7312 3394 8802 3453
rect 9140 3394 10630 3453
rect 10968 3394 12458 3453
rect 12796 3394 14286 3453
rect 14624 3394 16114 3453
rect 16452 3394 17942 3453
rect 18280 3394 19770 3453
rect 20108 3394 21598 3453
rect 22 3169 32 3322
rect 98 3169 108 3322
rect 214 3169 224 3322
rect 290 3169 300 3322
rect 406 3169 416 3322
rect 482 3169 492 3322
rect 598 3169 608 3322
rect 674 3169 684 3322
rect 790 3169 800 3322
rect 866 3169 876 3322
rect 982 3169 992 3322
rect 1058 3169 1068 3322
rect 1174 3169 1184 3322
rect 1250 3169 1260 3322
rect 1366 3169 1376 3322
rect 1442 3169 1452 3322
rect 1488 3109 1708 3356
rect 1850 3169 1860 3322
rect 1926 3169 1936 3322
rect 2042 3169 2052 3322
rect 2118 3169 2128 3322
rect 2234 3169 2244 3322
rect 2310 3169 2320 3322
rect 2426 3169 2436 3322
rect 2502 3169 2512 3322
rect 2618 3169 2628 3322
rect 2694 3169 2704 3322
rect 2810 3169 2820 3322
rect 2886 3169 2896 3322
rect 3002 3169 3012 3322
rect 3078 3169 3088 3322
rect 3194 3169 3204 3322
rect 3270 3169 3280 3322
rect 3316 3109 3536 3356
rect 3678 3169 3688 3322
rect 3754 3169 3764 3322
rect 3870 3169 3880 3322
rect 3946 3169 3956 3322
rect 4062 3169 4072 3322
rect 4138 3169 4148 3322
rect 4254 3169 4264 3322
rect 4330 3169 4340 3322
rect 4446 3169 4456 3322
rect 4522 3169 4532 3322
rect 4638 3169 4648 3322
rect 4714 3169 4724 3322
rect 4830 3169 4840 3322
rect 4906 3169 4916 3322
rect 5022 3169 5032 3322
rect 5098 3169 5108 3322
rect 5144 3109 5364 3356
rect 5506 3169 5516 3322
rect 5582 3169 5592 3322
rect 5698 3169 5708 3322
rect 5774 3169 5784 3322
rect 5890 3169 5900 3322
rect 5966 3169 5976 3322
rect 6082 3169 6092 3322
rect 6158 3169 6168 3322
rect 6274 3169 6284 3322
rect 6350 3169 6360 3322
rect 6466 3169 6476 3322
rect 6542 3169 6552 3322
rect 6658 3169 6668 3322
rect 6734 3169 6744 3322
rect 6850 3169 6860 3322
rect 6926 3169 6936 3322
rect 6972 3109 7192 3356
rect 7334 3169 7344 3322
rect 7410 3169 7420 3322
rect 7526 3169 7536 3322
rect 7602 3169 7612 3322
rect 7718 3169 7728 3322
rect 7794 3169 7804 3322
rect 7910 3169 7920 3322
rect 7986 3169 7996 3322
rect 8102 3169 8112 3322
rect 8178 3169 8188 3322
rect 8294 3169 8304 3322
rect 8370 3169 8380 3322
rect 8486 3169 8496 3322
rect 8562 3169 8572 3322
rect 8678 3169 8688 3322
rect 8754 3169 8764 3322
rect 8800 3109 9020 3356
rect 9162 3169 9172 3322
rect 9238 3169 9248 3322
rect 9354 3169 9364 3322
rect 9430 3169 9440 3322
rect 9546 3169 9556 3322
rect 9622 3169 9632 3322
rect 9738 3169 9748 3322
rect 9814 3169 9824 3322
rect 9930 3169 9940 3322
rect 10006 3169 10016 3322
rect 10122 3169 10132 3322
rect 10198 3169 10208 3322
rect 10314 3169 10324 3322
rect 10390 3169 10400 3322
rect 10506 3169 10516 3322
rect 10582 3169 10592 3322
rect 10628 3109 10848 3356
rect 10990 3169 11000 3322
rect 11066 3169 11076 3322
rect 11182 3169 11192 3322
rect 11258 3169 11268 3322
rect 11374 3169 11384 3322
rect 11450 3169 11460 3322
rect 11566 3169 11576 3322
rect 11642 3169 11652 3322
rect 11758 3169 11768 3322
rect 11834 3169 11844 3322
rect 11950 3169 11960 3322
rect 12026 3169 12036 3322
rect 12142 3169 12152 3322
rect 12218 3169 12228 3322
rect 12334 3169 12344 3322
rect 12410 3169 12420 3322
rect 12456 3109 12676 3356
rect 12818 3169 12828 3322
rect 12894 3169 12904 3322
rect 13010 3169 13020 3322
rect 13086 3169 13096 3322
rect 13202 3169 13212 3322
rect 13278 3169 13288 3322
rect 13394 3169 13404 3322
rect 13470 3169 13480 3322
rect 13586 3169 13596 3322
rect 13662 3169 13672 3322
rect 13778 3169 13788 3322
rect 13854 3169 13864 3322
rect 13970 3169 13980 3322
rect 14046 3169 14056 3322
rect 14162 3169 14172 3322
rect 14238 3169 14248 3322
rect 14284 3109 14504 3356
rect 14646 3169 14656 3322
rect 14722 3169 14732 3322
rect 14838 3169 14848 3322
rect 14914 3169 14924 3322
rect 15030 3169 15040 3322
rect 15106 3169 15116 3322
rect 15222 3169 15232 3322
rect 15298 3169 15308 3322
rect 15414 3169 15424 3322
rect 15490 3169 15500 3322
rect 15606 3169 15616 3322
rect 15682 3169 15692 3322
rect 15798 3169 15808 3322
rect 15874 3169 15884 3322
rect 15990 3169 16000 3322
rect 16066 3169 16076 3322
rect 16112 3109 16332 3356
rect 16474 3169 16484 3322
rect 16550 3169 16560 3322
rect 16666 3169 16676 3322
rect 16742 3169 16752 3322
rect 16858 3169 16868 3322
rect 16934 3169 16944 3322
rect 17050 3169 17060 3322
rect 17126 3169 17136 3322
rect 17242 3169 17252 3322
rect 17318 3169 17328 3322
rect 17434 3169 17444 3322
rect 17510 3169 17520 3322
rect 17626 3169 17636 3322
rect 17702 3169 17712 3322
rect 17818 3169 17828 3322
rect 17894 3169 17904 3322
rect 17940 3109 18160 3356
rect 18302 3169 18312 3322
rect 18378 3169 18388 3322
rect 18494 3169 18504 3322
rect 18570 3169 18580 3322
rect 18686 3169 18696 3322
rect 18762 3169 18772 3322
rect 18878 3169 18888 3322
rect 18954 3169 18964 3322
rect 19070 3169 19080 3322
rect 19146 3169 19156 3322
rect 19262 3169 19272 3322
rect 19338 3169 19348 3322
rect 19454 3169 19464 3322
rect 19530 3169 19540 3322
rect 19646 3169 19656 3322
rect 19722 3169 19732 3322
rect 19768 3109 19988 3356
rect 20130 3169 20140 3322
rect 20206 3169 20216 3322
rect 20322 3169 20332 3322
rect 20398 3169 20408 3322
rect 20514 3169 20524 3322
rect 20590 3169 20600 3322
rect 20706 3169 20716 3322
rect 20782 3169 20792 3322
rect 20898 3169 20908 3322
rect 20974 3169 20984 3322
rect 21090 3169 21100 3322
rect 21166 3169 21176 3322
rect 21282 3169 21292 3322
rect 21358 3169 21368 3322
rect 21474 3169 21484 3322
rect 21550 3169 21560 3322
rect 21596 3109 21816 3356
rect 118 2956 128 3109
rect 194 2956 204 3109
rect 310 2956 320 3109
rect 386 2956 396 3109
rect 502 2956 512 3109
rect 578 2956 588 3109
rect 694 2956 704 3109
rect 770 2956 780 3109
rect 886 2956 896 3109
rect 962 2956 972 3109
rect 1078 2956 1088 3109
rect 1154 2956 1164 3109
rect 1270 2956 1280 3109
rect 1346 2956 1356 3109
rect 1462 2956 1472 3109
rect 1528 2956 1708 3109
rect 1946 2956 1956 3109
rect 2022 2956 2032 3109
rect 2138 2956 2148 3109
rect 2214 2956 2224 3109
rect 2330 2956 2340 3109
rect 2406 2956 2416 3109
rect 2522 2956 2532 3109
rect 2598 2956 2608 3109
rect 2714 2956 2724 3109
rect 2790 2956 2800 3109
rect 2906 2956 2916 3109
rect 2982 2956 2992 3109
rect 3098 2956 3108 3109
rect 3174 2956 3184 3109
rect 3290 2956 3300 3109
rect 3356 2956 3536 3109
rect 3774 2956 3784 3109
rect 3850 2956 3860 3109
rect 3966 2956 3976 3109
rect 4042 2956 4052 3109
rect 4158 2956 4168 3109
rect 4234 2956 4244 3109
rect 4350 2956 4360 3109
rect 4426 2956 4436 3109
rect 4542 2956 4552 3109
rect 4618 2956 4628 3109
rect 4734 2956 4744 3109
rect 4810 2956 4820 3109
rect 4926 2956 4936 3109
rect 5002 2956 5012 3109
rect 5118 2956 5128 3109
rect 5184 2956 5364 3109
rect 5602 2956 5612 3109
rect 5678 2956 5688 3109
rect 5794 2956 5804 3109
rect 5870 2956 5880 3109
rect 5986 2956 5996 3109
rect 6062 2956 6072 3109
rect 6178 2956 6188 3109
rect 6254 2956 6264 3109
rect 6370 2956 6380 3109
rect 6446 2956 6456 3109
rect 6562 2956 6572 3109
rect 6638 2956 6648 3109
rect 6754 2956 6764 3109
rect 6830 2956 6840 3109
rect 6946 2956 6956 3109
rect 7012 2956 7192 3109
rect 7430 2956 7440 3109
rect 7506 2956 7516 3109
rect 7622 2956 7632 3109
rect 7698 2956 7708 3109
rect 7814 2956 7824 3109
rect 7890 2956 7900 3109
rect 8006 2956 8016 3109
rect 8082 2956 8092 3109
rect 8198 2956 8208 3109
rect 8274 2956 8284 3109
rect 8390 2956 8400 3109
rect 8466 2956 8476 3109
rect 8582 2956 8592 3109
rect 8658 2956 8668 3109
rect 8774 2956 8784 3109
rect 8840 2956 9020 3109
rect 9258 2956 9268 3109
rect 9334 2956 9344 3109
rect 9450 2956 9460 3109
rect 9526 2956 9536 3109
rect 9642 2956 9652 3109
rect 9718 2956 9728 3109
rect 9834 2956 9844 3109
rect 9910 2956 9920 3109
rect 10026 2956 10036 3109
rect 10102 2956 10112 3109
rect 10218 2956 10228 3109
rect 10294 2956 10304 3109
rect 10410 2956 10420 3109
rect 10486 2956 10496 3109
rect 10602 2956 10612 3109
rect 10668 2956 10848 3109
rect 11086 2956 11096 3109
rect 11162 2956 11172 3109
rect 11278 2956 11288 3109
rect 11354 2956 11364 3109
rect 11470 2956 11480 3109
rect 11546 2956 11556 3109
rect 11662 2956 11672 3109
rect 11738 2956 11748 3109
rect 11854 2956 11864 3109
rect 11930 2956 11940 3109
rect 12046 2956 12056 3109
rect 12122 2956 12132 3109
rect 12238 2956 12248 3109
rect 12314 2956 12324 3109
rect 12430 2956 12440 3109
rect 12496 2956 12676 3109
rect 12914 2956 12924 3109
rect 12990 2956 13000 3109
rect 13106 2956 13116 3109
rect 13182 2956 13192 3109
rect 13298 2956 13308 3109
rect 13374 2956 13384 3109
rect 13490 2956 13500 3109
rect 13566 2956 13576 3109
rect 13682 2956 13692 3109
rect 13758 2956 13768 3109
rect 13874 2956 13884 3109
rect 13950 2956 13960 3109
rect 14066 2956 14076 3109
rect 14142 2956 14152 3109
rect 14258 2956 14268 3109
rect 14324 2956 14504 3109
rect 14742 2956 14752 3109
rect 14818 2956 14828 3109
rect 14934 2956 14944 3109
rect 15010 2956 15020 3109
rect 15126 2956 15136 3109
rect 15202 2956 15212 3109
rect 15318 2956 15328 3109
rect 15394 2956 15404 3109
rect 15510 2956 15520 3109
rect 15586 2956 15596 3109
rect 15702 2956 15712 3109
rect 15778 2956 15788 3109
rect 15894 2956 15904 3109
rect 15970 2956 15980 3109
rect 16086 2956 16096 3109
rect 16152 2956 16332 3109
rect 16570 2956 16580 3109
rect 16646 2956 16656 3109
rect 16762 2956 16772 3109
rect 16838 2956 16848 3109
rect 16954 2956 16964 3109
rect 17030 2956 17040 3109
rect 17146 2956 17156 3109
rect 17222 2956 17232 3109
rect 17338 2956 17348 3109
rect 17414 2956 17424 3109
rect 17530 2956 17540 3109
rect 17606 2956 17616 3109
rect 17722 2956 17732 3109
rect 17798 2956 17808 3109
rect 17914 2956 17924 3109
rect 17980 2956 18160 3109
rect 18398 2956 18408 3109
rect 18474 2956 18484 3109
rect 18590 2956 18600 3109
rect 18666 2956 18676 3109
rect 18782 2956 18792 3109
rect 18858 2956 18868 3109
rect 18974 2956 18984 3109
rect 19050 2956 19060 3109
rect 19166 2956 19176 3109
rect 19242 2956 19252 3109
rect 19358 2956 19368 3109
rect 19434 2956 19444 3109
rect 19550 2956 19560 3109
rect 19626 2956 19636 3109
rect 19742 2956 19752 3109
rect 19808 2956 19988 3109
rect 20226 2956 20236 3109
rect 20302 2956 20312 3109
rect 20418 2956 20428 3109
rect 20494 2956 20504 3109
rect 20610 2956 20620 3109
rect 20686 2956 20696 3109
rect 20802 2956 20812 3109
rect 20878 2956 20888 3109
rect 20994 2956 21004 3109
rect 21070 2956 21080 3109
rect 21186 2956 21196 3109
rect 21262 2956 21272 3109
rect 21378 2956 21388 3109
rect 21454 2956 21464 3109
rect 21570 2956 21580 3109
rect 21636 2956 21816 3109
rect 0 2859 1490 2918
rect 1828 2859 3318 2918
rect 3656 2859 5146 2918
rect 5484 2859 6974 2918
rect 7312 2859 8802 2918
rect 9140 2859 10630 2918
rect 10968 2859 12458 2918
rect 12796 2859 14286 2918
rect 14624 2859 16114 2918
rect 16452 2859 17942 2918
rect 18280 2859 19770 2918
rect 20108 2859 21598 2918
rect 0 2680 1490 2739
rect 1828 2680 3318 2739
rect 3656 2680 5146 2739
rect 5484 2680 6974 2739
rect 7312 2680 8802 2739
rect 9140 2680 10630 2739
rect 10968 2680 12458 2739
rect 12796 2680 14286 2739
rect 14624 2680 16114 2739
rect 16452 2680 17942 2739
rect 18280 2680 19770 2739
rect 20108 2680 21598 2739
rect 22 2455 32 2608
rect 98 2455 108 2608
rect 214 2455 224 2608
rect 290 2455 300 2608
rect 406 2455 416 2608
rect 482 2455 492 2608
rect 598 2455 608 2608
rect 674 2455 684 2608
rect 790 2455 800 2608
rect 866 2455 876 2608
rect 982 2455 992 2608
rect 1058 2455 1068 2608
rect 1174 2455 1184 2608
rect 1250 2455 1260 2608
rect 1366 2455 1376 2608
rect 1442 2455 1452 2608
rect 1488 2395 1708 2642
rect 1850 2455 1860 2608
rect 1926 2455 1936 2608
rect 2042 2455 2052 2608
rect 2118 2455 2128 2608
rect 2234 2455 2244 2608
rect 2310 2455 2320 2608
rect 2426 2455 2436 2608
rect 2502 2455 2512 2608
rect 2618 2455 2628 2608
rect 2694 2455 2704 2608
rect 2810 2455 2820 2608
rect 2886 2455 2896 2608
rect 3002 2455 3012 2608
rect 3078 2455 3088 2608
rect 3194 2455 3204 2608
rect 3270 2455 3280 2608
rect 3316 2395 3536 2642
rect 3678 2455 3688 2608
rect 3754 2455 3764 2608
rect 3870 2455 3880 2608
rect 3946 2455 3956 2608
rect 4062 2455 4072 2608
rect 4138 2455 4148 2608
rect 4254 2455 4264 2608
rect 4330 2455 4340 2608
rect 4446 2455 4456 2608
rect 4522 2455 4532 2608
rect 4638 2455 4648 2608
rect 4714 2455 4724 2608
rect 4830 2455 4840 2608
rect 4906 2455 4916 2608
rect 5022 2455 5032 2608
rect 5098 2455 5108 2608
rect 5144 2395 5364 2642
rect 5506 2455 5516 2608
rect 5582 2455 5592 2608
rect 5698 2455 5708 2608
rect 5774 2455 5784 2608
rect 5890 2455 5900 2608
rect 5966 2455 5976 2608
rect 6082 2455 6092 2608
rect 6158 2455 6168 2608
rect 6274 2455 6284 2608
rect 6350 2455 6360 2608
rect 6466 2455 6476 2608
rect 6542 2455 6552 2608
rect 6658 2455 6668 2608
rect 6734 2455 6744 2608
rect 6850 2455 6860 2608
rect 6926 2455 6936 2608
rect 6972 2395 7192 2642
rect 7334 2455 7344 2608
rect 7410 2455 7420 2608
rect 7526 2455 7536 2608
rect 7602 2455 7612 2608
rect 7718 2455 7728 2608
rect 7794 2455 7804 2608
rect 7910 2455 7920 2608
rect 7986 2455 7996 2608
rect 8102 2455 8112 2608
rect 8178 2455 8188 2608
rect 8294 2455 8304 2608
rect 8370 2455 8380 2608
rect 8486 2455 8496 2608
rect 8562 2455 8572 2608
rect 8678 2455 8688 2608
rect 8754 2455 8764 2608
rect 8800 2395 9020 2642
rect 9162 2455 9172 2608
rect 9238 2455 9248 2608
rect 9354 2455 9364 2608
rect 9430 2455 9440 2608
rect 9546 2455 9556 2608
rect 9622 2455 9632 2608
rect 9738 2455 9748 2608
rect 9814 2455 9824 2608
rect 9930 2455 9940 2608
rect 10006 2455 10016 2608
rect 10122 2455 10132 2608
rect 10198 2455 10208 2608
rect 10314 2455 10324 2608
rect 10390 2455 10400 2608
rect 10506 2455 10516 2608
rect 10582 2455 10592 2608
rect 10628 2395 10848 2642
rect 10990 2455 11000 2608
rect 11066 2455 11076 2608
rect 11182 2455 11192 2608
rect 11258 2455 11268 2608
rect 11374 2455 11384 2608
rect 11450 2455 11460 2608
rect 11566 2455 11576 2608
rect 11642 2455 11652 2608
rect 11758 2455 11768 2608
rect 11834 2455 11844 2608
rect 11950 2455 11960 2608
rect 12026 2455 12036 2608
rect 12142 2455 12152 2608
rect 12218 2455 12228 2608
rect 12334 2455 12344 2608
rect 12410 2455 12420 2608
rect 12456 2395 12676 2642
rect 12818 2455 12828 2608
rect 12894 2455 12904 2608
rect 13010 2455 13020 2608
rect 13086 2455 13096 2608
rect 13202 2455 13212 2608
rect 13278 2455 13288 2608
rect 13394 2455 13404 2608
rect 13470 2455 13480 2608
rect 13586 2455 13596 2608
rect 13662 2455 13672 2608
rect 13778 2455 13788 2608
rect 13854 2455 13864 2608
rect 13970 2455 13980 2608
rect 14046 2455 14056 2608
rect 14162 2455 14172 2608
rect 14238 2455 14248 2608
rect 14284 2395 14504 2642
rect 14646 2455 14656 2608
rect 14722 2455 14732 2608
rect 14838 2455 14848 2608
rect 14914 2455 14924 2608
rect 15030 2455 15040 2608
rect 15106 2455 15116 2608
rect 15222 2455 15232 2608
rect 15298 2455 15308 2608
rect 15414 2455 15424 2608
rect 15490 2455 15500 2608
rect 15606 2455 15616 2608
rect 15682 2455 15692 2608
rect 15798 2455 15808 2608
rect 15874 2455 15884 2608
rect 15990 2455 16000 2608
rect 16066 2455 16076 2608
rect 16112 2395 16332 2642
rect 16474 2455 16484 2608
rect 16550 2455 16560 2608
rect 16666 2455 16676 2608
rect 16742 2455 16752 2608
rect 16858 2455 16868 2608
rect 16934 2455 16944 2608
rect 17050 2455 17060 2608
rect 17126 2455 17136 2608
rect 17242 2455 17252 2608
rect 17318 2455 17328 2608
rect 17434 2455 17444 2608
rect 17510 2455 17520 2608
rect 17626 2455 17636 2608
rect 17702 2455 17712 2608
rect 17818 2455 17828 2608
rect 17894 2455 17904 2608
rect 17940 2395 18160 2642
rect 18302 2455 18312 2608
rect 18378 2455 18388 2608
rect 18494 2455 18504 2608
rect 18570 2455 18580 2608
rect 18686 2455 18696 2608
rect 18762 2455 18772 2608
rect 18878 2455 18888 2608
rect 18954 2455 18964 2608
rect 19070 2455 19080 2608
rect 19146 2455 19156 2608
rect 19262 2455 19272 2608
rect 19338 2455 19348 2608
rect 19454 2455 19464 2608
rect 19530 2455 19540 2608
rect 19646 2455 19656 2608
rect 19722 2455 19732 2608
rect 19768 2395 19988 2642
rect 20130 2455 20140 2608
rect 20206 2455 20216 2608
rect 20322 2455 20332 2608
rect 20398 2455 20408 2608
rect 20514 2455 20524 2608
rect 20590 2455 20600 2608
rect 20706 2455 20716 2608
rect 20782 2455 20792 2608
rect 20898 2455 20908 2608
rect 20974 2455 20984 2608
rect 21090 2455 21100 2608
rect 21166 2455 21176 2608
rect 21282 2455 21292 2608
rect 21358 2455 21368 2608
rect 21474 2455 21484 2608
rect 21550 2455 21560 2608
rect 21596 2395 21816 2642
rect 118 2242 128 2395
rect 194 2242 204 2395
rect 310 2242 320 2395
rect 386 2242 396 2395
rect 502 2242 512 2395
rect 578 2242 588 2395
rect 694 2242 704 2395
rect 770 2242 780 2395
rect 886 2242 896 2395
rect 962 2242 972 2395
rect 1078 2242 1088 2395
rect 1154 2242 1164 2395
rect 1270 2242 1280 2395
rect 1346 2242 1356 2395
rect 1462 2242 1472 2395
rect 1528 2242 1708 2395
rect 1946 2242 1956 2395
rect 2022 2242 2032 2395
rect 2138 2242 2148 2395
rect 2214 2242 2224 2395
rect 2330 2242 2340 2395
rect 2406 2242 2416 2395
rect 2522 2242 2532 2395
rect 2598 2242 2608 2395
rect 2714 2242 2724 2395
rect 2790 2242 2800 2395
rect 2906 2242 2916 2395
rect 2982 2242 2992 2395
rect 3098 2242 3108 2395
rect 3174 2242 3184 2395
rect 3290 2242 3300 2395
rect 3356 2242 3536 2395
rect 3774 2242 3784 2395
rect 3850 2242 3860 2395
rect 3966 2242 3976 2395
rect 4042 2242 4052 2395
rect 4158 2242 4168 2395
rect 4234 2242 4244 2395
rect 4350 2242 4360 2395
rect 4426 2242 4436 2395
rect 4542 2242 4552 2395
rect 4618 2242 4628 2395
rect 4734 2242 4744 2395
rect 4810 2242 4820 2395
rect 4926 2242 4936 2395
rect 5002 2242 5012 2395
rect 5118 2242 5128 2395
rect 5184 2242 5364 2395
rect 5602 2242 5612 2395
rect 5678 2242 5688 2395
rect 5794 2242 5804 2395
rect 5870 2242 5880 2395
rect 5986 2242 5996 2395
rect 6062 2242 6072 2395
rect 6178 2242 6188 2395
rect 6254 2242 6264 2395
rect 6370 2242 6380 2395
rect 6446 2242 6456 2395
rect 6562 2242 6572 2395
rect 6638 2242 6648 2395
rect 6754 2242 6764 2395
rect 6830 2242 6840 2395
rect 6946 2242 6956 2395
rect 7012 2242 7192 2395
rect 7430 2242 7440 2395
rect 7506 2242 7516 2395
rect 7622 2242 7632 2395
rect 7698 2242 7708 2395
rect 7814 2242 7824 2395
rect 7890 2242 7900 2395
rect 8006 2242 8016 2395
rect 8082 2242 8092 2395
rect 8198 2242 8208 2395
rect 8274 2242 8284 2395
rect 8390 2242 8400 2395
rect 8466 2242 8476 2395
rect 8582 2242 8592 2395
rect 8658 2242 8668 2395
rect 8774 2242 8784 2395
rect 8840 2242 9020 2395
rect 9258 2242 9268 2395
rect 9334 2242 9344 2395
rect 9450 2242 9460 2395
rect 9526 2242 9536 2395
rect 9642 2242 9652 2395
rect 9718 2242 9728 2395
rect 9834 2242 9844 2395
rect 9910 2242 9920 2395
rect 10026 2242 10036 2395
rect 10102 2242 10112 2395
rect 10218 2242 10228 2395
rect 10294 2242 10304 2395
rect 10410 2242 10420 2395
rect 10486 2242 10496 2395
rect 10602 2242 10612 2395
rect 10668 2242 10848 2395
rect 11086 2242 11096 2395
rect 11162 2242 11172 2395
rect 11278 2242 11288 2395
rect 11354 2242 11364 2395
rect 11470 2242 11480 2395
rect 11546 2242 11556 2395
rect 11662 2242 11672 2395
rect 11738 2242 11748 2395
rect 11854 2242 11864 2395
rect 11930 2242 11940 2395
rect 12046 2242 12056 2395
rect 12122 2242 12132 2395
rect 12238 2242 12248 2395
rect 12314 2242 12324 2395
rect 12430 2242 12440 2395
rect 12496 2242 12676 2395
rect 12914 2242 12924 2395
rect 12990 2242 13000 2395
rect 13106 2242 13116 2395
rect 13182 2242 13192 2395
rect 13298 2242 13308 2395
rect 13374 2242 13384 2395
rect 13490 2242 13500 2395
rect 13566 2242 13576 2395
rect 13682 2242 13692 2395
rect 13758 2242 13768 2395
rect 13874 2242 13884 2395
rect 13950 2242 13960 2395
rect 14066 2242 14076 2395
rect 14142 2242 14152 2395
rect 14258 2242 14268 2395
rect 14324 2242 14504 2395
rect 14742 2242 14752 2395
rect 14818 2242 14828 2395
rect 14934 2242 14944 2395
rect 15010 2242 15020 2395
rect 15126 2242 15136 2395
rect 15202 2242 15212 2395
rect 15318 2242 15328 2395
rect 15394 2242 15404 2395
rect 15510 2242 15520 2395
rect 15586 2242 15596 2395
rect 15702 2242 15712 2395
rect 15778 2242 15788 2395
rect 15894 2242 15904 2395
rect 15970 2242 15980 2395
rect 16086 2242 16096 2395
rect 16152 2242 16332 2395
rect 16570 2242 16580 2395
rect 16646 2242 16656 2395
rect 16762 2242 16772 2395
rect 16838 2242 16848 2395
rect 16954 2242 16964 2395
rect 17030 2242 17040 2395
rect 17146 2242 17156 2395
rect 17222 2242 17232 2395
rect 17338 2242 17348 2395
rect 17414 2242 17424 2395
rect 17530 2242 17540 2395
rect 17606 2242 17616 2395
rect 17722 2242 17732 2395
rect 17798 2242 17808 2395
rect 17914 2242 17924 2395
rect 17980 2242 18160 2395
rect 18398 2242 18408 2395
rect 18474 2242 18484 2395
rect 18590 2242 18600 2395
rect 18666 2242 18676 2395
rect 18782 2242 18792 2395
rect 18858 2242 18868 2395
rect 18974 2242 18984 2395
rect 19050 2242 19060 2395
rect 19166 2242 19176 2395
rect 19242 2242 19252 2395
rect 19358 2242 19368 2395
rect 19434 2242 19444 2395
rect 19550 2242 19560 2395
rect 19626 2242 19636 2395
rect 19742 2242 19752 2395
rect 19808 2242 19988 2395
rect 20226 2242 20236 2395
rect 20302 2242 20312 2395
rect 20418 2242 20428 2395
rect 20494 2242 20504 2395
rect 20610 2242 20620 2395
rect 20686 2242 20696 2395
rect 20802 2242 20812 2395
rect 20878 2242 20888 2395
rect 20994 2242 21004 2395
rect 21070 2242 21080 2395
rect 21186 2242 21196 2395
rect 21262 2242 21272 2395
rect 21378 2242 21388 2395
rect 21454 2242 21464 2395
rect 21570 2242 21580 2395
rect 21636 2242 21816 2395
rect 0 2145 1490 2204
rect 1828 2145 3318 2204
rect 3656 2145 5146 2204
rect 5484 2145 6974 2204
rect 7312 2145 8802 2204
rect 9140 2145 10630 2204
rect 10968 2145 12458 2204
rect 12796 2145 14286 2204
rect 14624 2145 16114 2204
rect 16452 2145 17942 2204
rect 18280 2145 19770 2204
rect 20108 2145 21598 2204
rect 0 1966 1490 2025
rect 1828 1966 3318 2025
rect 3656 1966 5146 2025
rect 5484 1966 6974 2025
rect 7312 1966 8802 2025
rect 9140 1966 10630 2025
rect 10968 1966 12458 2025
rect 12796 1966 14286 2025
rect 14624 1966 16114 2025
rect 16452 1966 17942 2025
rect 18280 1966 19770 2025
rect 20108 1966 21598 2025
rect 22 1741 32 1894
rect 98 1741 108 1894
rect 214 1741 224 1894
rect 290 1741 300 1894
rect 406 1741 416 1894
rect 482 1741 492 1894
rect 598 1741 608 1894
rect 674 1741 684 1894
rect 790 1741 800 1894
rect 866 1741 876 1894
rect 982 1741 992 1894
rect 1058 1741 1068 1894
rect 1174 1741 1184 1894
rect 1250 1741 1260 1894
rect 1366 1741 1376 1894
rect 1442 1741 1452 1894
rect 1488 1681 1708 1928
rect 1850 1741 1860 1894
rect 1926 1741 1936 1894
rect 2042 1741 2052 1894
rect 2118 1741 2128 1894
rect 2234 1741 2244 1894
rect 2310 1741 2320 1894
rect 2426 1741 2436 1894
rect 2502 1741 2512 1894
rect 2618 1741 2628 1894
rect 2694 1741 2704 1894
rect 2810 1741 2820 1894
rect 2886 1741 2896 1894
rect 3002 1741 3012 1894
rect 3078 1741 3088 1894
rect 3194 1741 3204 1894
rect 3270 1741 3280 1894
rect 3316 1681 3536 1928
rect 3678 1741 3688 1894
rect 3754 1741 3764 1894
rect 3870 1741 3880 1894
rect 3946 1741 3956 1894
rect 4062 1741 4072 1894
rect 4138 1741 4148 1894
rect 4254 1741 4264 1894
rect 4330 1741 4340 1894
rect 4446 1741 4456 1894
rect 4522 1741 4532 1894
rect 4638 1741 4648 1894
rect 4714 1741 4724 1894
rect 4830 1741 4840 1894
rect 4906 1741 4916 1894
rect 5022 1741 5032 1894
rect 5098 1741 5108 1894
rect 5144 1681 5364 1928
rect 5506 1741 5516 1894
rect 5582 1741 5592 1894
rect 5698 1741 5708 1894
rect 5774 1741 5784 1894
rect 5890 1741 5900 1894
rect 5966 1741 5976 1894
rect 6082 1741 6092 1894
rect 6158 1741 6168 1894
rect 6274 1741 6284 1894
rect 6350 1741 6360 1894
rect 6466 1741 6476 1894
rect 6542 1741 6552 1894
rect 6658 1741 6668 1894
rect 6734 1741 6744 1894
rect 6850 1741 6860 1894
rect 6926 1741 6936 1894
rect 6972 1681 7192 1928
rect 7334 1741 7344 1894
rect 7410 1741 7420 1894
rect 7526 1741 7536 1894
rect 7602 1741 7612 1894
rect 7718 1741 7728 1894
rect 7794 1741 7804 1894
rect 7910 1741 7920 1894
rect 7986 1741 7996 1894
rect 8102 1741 8112 1894
rect 8178 1741 8188 1894
rect 8294 1741 8304 1894
rect 8370 1741 8380 1894
rect 8486 1741 8496 1894
rect 8562 1741 8572 1894
rect 8678 1741 8688 1894
rect 8754 1741 8764 1894
rect 8800 1681 9020 1928
rect 9162 1741 9172 1894
rect 9238 1741 9248 1894
rect 9354 1741 9364 1894
rect 9430 1741 9440 1894
rect 9546 1741 9556 1894
rect 9622 1741 9632 1894
rect 9738 1741 9748 1894
rect 9814 1741 9824 1894
rect 9930 1741 9940 1894
rect 10006 1741 10016 1894
rect 10122 1741 10132 1894
rect 10198 1741 10208 1894
rect 10314 1741 10324 1894
rect 10390 1741 10400 1894
rect 10506 1741 10516 1894
rect 10582 1741 10592 1894
rect 10628 1681 10848 1928
rect 10990 1741 11000 1894
rect 11066 1741 11076 1894
rect 11182 1741 11192 1894
rect 11258 1741 11268 1894
rect 11374 1741 11384 1894
rect 11450 1741 11460 1894
rect 11566 1741 11576 1894
rect 11642 1741 11652 1894
rect 11758 1741 11768 1894
rect 11834 1741 11844 1894
rect 11950 1741 11960 1894
rect 12026 1741 12036 1894
rect 12142 1741 12152 1894
rect 12218 1741 12228 1894
rect 12334 1741 12344 1894
rect 12410 1741 12420 1894
rect 12456 1681 12676 1928
rect 12818 1741 12828 1894
rect 12894 1741 12904 1894
rect 13010 1741 13020 1894
rect 13086 1741 13096 1894
rect 13202 1741 13212 1894
rect 13278 1741 13288 1894
rect 13394 1741 13404 1894
rect 13470 1741 13480 1894
rect 13586 1741 13596 1894
rect 13662 1741 13672 1894
rect 13778 1741 13788 1894
rect 13854 1741 13864 1894
rect 13970 1741 13980 1894
rect 14046 1741 14056 1894
rect 14162 1741 14172 1894
rect 14238 1741 14248 1894
rect 14284 1681 14504 1928
rect 14646 1741 14656 1894
rect 14722 1741 14732 1894
rect 14838 1741 14848 1894
rect 14914 1741 14924 1894
rect 15030 1741 15040 1894
rect 15106 1741 15116 1894
rect 15222 1741 15232 1894
rect 15298 1741 15308 1894
rect 15414 1741 15424 1894
rect 15490 1741 15500 1894
rect 15606 1741 15616 1894
rect 15682 1741 15692 1894
rect 15798 1741 15808 1894
rect 15874 1741 15884 1894
rect 15990 1741 16000 1894
rect 16066 1741 16076 1894
rect 16112 1681 16332 1928
rect 16474 1741 16484 1894
rect 16550 1741 16560 1894
rect 16666 1741 16676 1894
rect 16742 1741 16752 1894
rect 16858 1741 16868 1894
rect 16934 1741 16944 1894
rect 17050 1741 17060 1894
rect 17126 1741 17136 1894
rect 17242 1741 17252 1894
rect 17318 1741 17328 1894
rect 17434 1741 17444 1894
rect 17510 1741 17520 1894
rect 17626 1741 17636 1894
rect 17702 1741 17712 1894
rect 17818 1741 17828 1894
rect 17894 1741 17904 1894
rect 17940 1681 18160 1928
rect 18302 1741 18312 1894
rect 18378 1741 18388 1894
rect 18494 1741 18504 1894
rect 18570 1741 18580 1894
rect 18686 1741 18696 1894
rect 18762 1741 18772 1894
rect 18878 1741 18888 1894
rect 18954 1741 18964 1894
rect 19070 1741 19080 1894
rect 19146 1741 19156 1894
rect 19262 1741 19272 1894
rect 19338 1741 19348 1894
rect 19454 1741 19464 1894
rect 19530 1741 19540 1894
rect 19646 1741 19656 1894
rect 19722 1741 19732 1894
rect 19768 1681 19988 1928
rect 20130 1741 20140 1894
rect 20206 1741 20216 1894
rect 20322 1741 20332 1894
rect 20398 1741 20408 1894
rect 20514 1741 20524 1894
rect 20590 1741 20600 1894
rect 20706 1741 20716 1894
rect 20782 1741 20792 1894
rect 20898 1741 20908 1894
rect 20974 1741 20984 1894
rect 21090 1741 21100 1894
rect 21166 1741 21176 1894
rect 21282 1741 21292 1894
rect 21358 1741 21368 1894
rect 21474 1741 21484 1894
rect 21550 1741 21560 1894
rect 21596 1681 21816 1928
rect 118 1528 128 1681
rect 194 1528 204 1681
rect 310 1528 320 1681
rect 386 1528 396 1681
rect 502 1528 512 1681
rect 578 1528 588 1681
rect 694 1528 704 1681
rect 770 1528 780 1681
rect 886 1528 896 1681
rect 962 1528 972 1681
rect 1078 1528 1088 1681
rect 1154 1528 1164 1681
rect 1270 1528 1280 1681
rect 1346 1528 1356 1681
rect 1462 1528 1472 1681
rect 1528 1528 1708 1681
rect 1946 1528 1956 1681
rect 2022 1528 2032 1681
rect 2138 1528 2148 1681
rect 2214 1528 2224 1681
rect 2330 1528 2340 1681
rect 2406 1528 2416 1681
rect 2522 1528 2532 1681
rect 2598 1528 2608 1681
rect 2714 1528 2724 1681
rect 2790 1528 2800 1681
rect 2906 1528 2916 1681
rect 2982 1528 2992 1681
rect 3098 1528 3108 1681
rect 3174 1528 3184 1681
rect 3290 1528 3300 1681
rect 3356 1528 3536 1681
rect 3774 1528 3784 1681
rect 3850 1528 3860 1681
rect 3966 1528 3976 1681
rect 4042 1528 4052 1681
rect 4158 1528 4168 1681
rect 4234 1528 4244 1681
rect 4350 1528 4360 1681
rect 4426 1528 4436 1681
rect 4542 1528 4552 1681
rect 4618 1528 4628 1681
rect 4734 1528 4744 1681
rect 4810 1528 4820 1681
rect 4926 1528 4936 1681
rect 5002 1528 5012 1681
rect 5118 1528 5128 1681
rect 5184 1528 5364 1681
rect 5602 1528 5612 1681
rect 5678 1528 5688 1681
rect 5794 1528 5804 1681
rect 5870 1528 5880 1681
rect 5986 1528 5996 1681
rect 6062 1528 6072 1681
rect 6178 1528 6188 1681
rect 6254 1528 6264 1681
rect 6370 1528 6380 1681
rect 6446 1528 6456 1681
rect 6562 1528 6572 1681
rect 6638 1528 6648 1681
rect 6754 1528 6764 1681
rect 6830 1528 6840 1681
rect 6946 1528 6956 1681
rect 7012 1528 7192 1681
rect 7430 1528 7440 1681
rect 7506 1528 7516 1681
rect 7622 1528 7632 1681
rect 7698 1528 7708 1681
rect 7814 1528 7824 1681
rect 7890 1528 7900 1681
rect 8006 1528 8016 1681
rect 8082 1528 8092 1681
rect 8198 1528 8208 1681
rect 8274 1528 8284 1681
rect 8390 1528 8400 1681
rect 8466 1528 8476 1681
rect 8582 1528 8592 1681
rect 8658 1528 8668 1681
rect 8774 1528 8784 1681
rect 8840 1528 9020 1681
rect 9258 1528 9268 1681
rect 9334 1528 9344 1681
rect 9450 1528 9460 1681
rect 9526 1528 9536 1681
rect 9642 1528 9652 1681
rect 9718 1528 9728 1681
rect 9834 1528 9844 1681
rect 9910 1528 9920 1681
rect 10026 1528 10036 1681
rect 10102 1528 10112 1681
rect 10218 1528 10228 1681
rect 10294 1528 10304 1681
rect 10410 1528 10420 1681
rect 10486 1528 10496 1681
rect 10602 1528 10612 1681
rect 10668 1528 10848 1681
rect 11086 1528 11096 1681
rect 11162 1528 11172 1681
rect 11278 1528 11288 1681
rect 11354 1528 11364 1681
rect 11470 1528 11480 1681
rect 11546 1528 11556 1681
rect 11662 1528 11672 1681
rect 11738 1528 11748 1681
rect 11854 1528 11864 1681
rect 11930 1528 11940 1681
rect 12046 1528 12056 1681
rect 12122 1528 12132 1681
rect 12238 1528 12248 1681
rect 12314 1528 12324 1681
rect 12430 1528 12440 1681
rect 12496 1528 12676 1681
rect 12914 1528 12924 1681
rect 12990 1528 13000 1681
rect 13106 1528 13116 1681
rect 13182 1528 13192 1681
rect 13298 1528 13308 1681
rect 13374 1528 13384 1681
rect 13490 1528 13500 1681
rect 13566 1528 13576 1681
rect 13682 1528 13692 1681
rect 13758 1528 13768 1681
rect 13874 1528 13884 1681
rect 13950 1528 13960 1681
rect 14066 1528 14076 1681
rect 14142 1528 14152 1681
rect 14258 1528 14268 1681
rect 14324 1528 14504 1681
rect 14742 1528 14752 1681
rect 14818 1528 14828 1681
rect 14934 1528 14944 1681
rect 15010 1528 15020 1681
rect 15126 1528 15136 1681
rect 15202 1528 15212 1681
rect 15318 1528 15328 1681
rect 15394 1528 15404 1681
rect 15510 1528 15520 1681
rect 15586 1528 15596 1681
rect 15702 1528 15712 1681
rect 15778 1528 15788 1681
rect 15894 1528 15904 1681
rect 15970 1528 15980 1681
rect 16086 1528 16096 1681
rect 16152 1528 16332 1681
rect 16570 1528 16580 1681
rect 16646 1528 16656 1681
rect 16762 1528 16772 1681
rect 16838 1528 16848 1681
rect 16954 1528 16964 1681
rect 17030 1528 17040 1681
rect 17146 1528 17156 1681
rect 17222 1528 17232 1681
rect 17338 1528 17348 1681
rect 17414 1528 17424 1681
rect 17530 1528 17540 1681
rect 17606 1528 17616 1681
rect 17722 1528 17732 1681
rect 17798 1528 17808 1681
rect 17914 1528 17924 1681
rect 17980 1528 18160 1681
rect 18398 1528 18408 1681
rect 18474 1528 18484 1681
rect 18590 1528 18600 1681
rect 18666 1528 18676 1681
rect 18782 1528 18792 1681
rect 18858 1528 18868 1681
rect 18974 1528 18984 1681
rect 19050 1528 19060 1681
rect 19166 1528 19176 1681
rect 19242 1528 19252 1681
rect 19358 1528 19368 1681
rect 19434 1528 19444 1681
rect 19550 1528 19560 1681
rect 19626 1528 19636 1681
rect 19742 1528 19752 1681
rect 19808 1528 19988 1681
rect 20226 1528 20236 1681
rect 20302 1528 20312 1681
rect 20418 1528 20428 1681
rect 20494 1528 20504 1681
rect 20610 1528 20620 1681
rect 20686 1528 20696 1681
rect 20802 1528 20812 1681
rect 20878 1528 20888 1681
rect 20994 1528 21004 1681
rect 21070 1528 21080 1681
rect 21186 1528 21196 1681
rect 21262 1528 21272 1681
rect 21378 1528 21388 1681
rect 21454 1528 21464 1681
rect 21570 1528 21580 1681
rect 21636 1528 21816 1681
rect 0 1431 1490 1490
rect 1828 1431 3318 1490
rect 3656 1431 5146 1490
rect 5484 1431 6974 1490
rect 7312 1431 8802 1490
rect 9140 1431 10630 1490
rect 10968 1431 12458 1490
rect 12796 1431 14286 1490
rect 14624 1431 16114 1490
rect 16452 1431 17942 1490
rect 18280 1431 19770 1490
rect 20108 1431 21598 1490
rect 0 1252 1490 1311
rect 1828 1252 3318 1311
rect 3656 1252 5146 1311
rect 5484 1252 6974 1311
rect 7312 1252 8802 1311
rect 9140 1252 10630 1311
rect 10968 1252 12458 1311
rect 12796 1252 14286 1311
rect 14624 1252 16114 1311
rect 16452 1252 17942 1311
rect 18280 1252 19770 1311
rect 20108 1252 21598 1311
rect 22 1027 32 1180
rect 98 1027 108 1180
rect 214 1027 224 1180
rect 290 1027 300 1180
rect 406 1027 416 1180
rect 482 1027 492 1180
rect 598 1027 608 1180
rect 674 1027 684 1180
rect 790 1027 800 1180
rect 866 1027 876 1180
rect 982 1027 992 1180
rect 1058 1027 1068 1180
rect 1174 1027 1184 1180
rect 1250 1027 1260 1180
rect 1366 1027 1376 1180
rect 1442 1027 1452 1180
rect 1488 967 1708 1214
rect 1850 1027 1860 1180
rect 1926 1027 1936 1180
rect 2042 1027 2052 1180
rect 2118 1027 2128 1180
rect 2234 1027 2244 1180
rect 2310 1027 2320 1180
rect 2426 1027 2436 1180
rect 2502 1027 2512 1180
rect 2618 1027 2628 1180
rect 2694 1027 2704 1180
rect 2810 1027 2820 1180
rect 2886 1027 2896 1180
rect 3002 1027 3012 1180
rect 3078 1027 3088 1180
rect 3194 1027 3204 1180
rect 3270 1027 3280 1180
rect 3316 967 3536 1214
rect 3678 1027 3688 1180
rect 3754 1027 3764 1180
rect 3870 1027 3880 1180
rect 3946 1027 3956 1180
rect 4062 1027 4072 1180
rect 4138 1027 4148 1180
rect 4254 1027 4264 1180
rect 4330 1027 4340 1180
rect 4446 1027 4456 1180
rect 4522 1027 4532 1180
rect 4638 1027 4648 1180
rect 4714 1027 4724 1180
rect 4830 1027 4840 1180
rect 4906 1027 4916 1180
rect 5022 1027 5032 1180
rect 5098 1027 5108 1180
rect 5144 967 5364 1214
rect 5506 1027 5516 1180
rect 5582 1027 5592 1180
rect 5698 1027 5708 1180
rect 5774 1027 5784 1180
rect 5890 1027 5900 1180
rect 5966 1027 5976 1180
rect 6082 1027 6092 1180
rect 6158 1027 6168 1180
rect 6274 1027 6284 1180
rect 6350 1027 6360 1180
rect 6466 1027 6476 1180
rect 6542 1027 6552 1180
rect 6658 1027 6668 1180
rect 6734 1027 6744 1180
rect 6850 1027 6860 1180
rect 6926 1027 6936 1180
rect 6972 967 7192 1214
rect 7334 1027 7344 1180
rect 7410 1027 7420 1180
rect 7526 1027 7536 1180
rect 7602 1027 7612 1180
rect 7718 1027 7728 1180
rect 7794 1027 7804 1180
rect 7910 1027 7920 1180
rect 7986 1027 7996 1180
rect 8102 1027 8112 1180
rect 8178 1027 8188 1180
rect 8294 1027 8304 1180
rect 8370 1027 8380 1180
rect 8486 1027 8496 1180
rect 8562 1027 8572 1180
rect 8678 1027 8688 1180
rect 8754 1027 8764 1180
rect 8800 967 9020 1214
rect 9162 1027 9172 1180
rect 9238 1027 9248 1180
rect 9354 1027 9364 1180
rect 9430 1027 9440 1180
rect 9546 1027 9556 1180
rect 9622 1027 9632 1180
rect 9738 1027 9748 1180
rect 9814 1027 9824 1180
rect 9930 1027 9940 1180
rect 10006 1027 10016 1180
rect 10122 1027 10132 1180
rect 10198 1027 10208 1180
rect 10314 1027 10324 1180
rect 10390 1027 10400 1180
rect 10506 1027 10516 1180
rect 10582 1027 10592 1180
rect 10628 967 10848 1214
rect 10990 1027 11000 1180
rect 11066 1027 11076 1180
rect 11182 1027 11192 1180
rect 11258 1027 11268 1180
rect 11374 1027 11384 1180
rect 11450 1027 11460 1180
rect 11566 1027 11576 1180
rect 11642 1027 11652 1180
rect 11758 1027 11768 1180
rect 11834 1027 11844 1180
rect 11950 1027 11960 1180
rect 12026 1027 12036 1180
rect 12142 1027 12152 1180
rect 12218 1027 12228 1180
rect 12334 1027 12344 1180
rect 12410 1027 12420 1180
rect 12456 967 12676 1214
rect 12818 1027 12828 1180
rect 12894 1027 12904 1180
rect 13010 1027 13020 1180
rect 13086 1027 13096 1180
rect 13202 1027 13212 1180
rect 13278 1027 13288 1180
rect 13394 1027 13404 1180
rect 13470 1027 13480 1180
rect 13586 1027 13596 1180
rect 13662 1027 13672 1180
rect 13778 1027 13788 1180
rect 13854 1027 13864 1180
rect 13970 1027 13980 1180
rect 14046 1027 14056 1180
rect 14162 1027 14172 1180
rect 14238 1027 14248 1180
rect 14284 967 14504 1214
rect 14646 1027 14656 1180
rect 14722 1027 14732 1180
rect 14838 1027 14848 1180
rect 14914 1027 14924 1180
rect 15030 1027 15040 1180
rect 15106 1027 15116 1180
rect 15222 1027 15232 1180
rect 15298 1027 15308 1180
rect 15414 1027 15424 1180
rect 15490 1027 15500 1180
rect 15606 1027 15616 1180
rect 15682 1027 15692 1180
rect 15798 1027 15808 1180
rect 15874 1027 15884 1180
rect 15990 1027 16000 1180
rect 16066 1027 16076 1180
rect 16112 967 16332 1214
rect 16474 1027 16484 1180
rect 16550 1027 16560 1180
rect 16666 1027 16676 1180
rect 16742 1027 16752 1180
rect 16858 1027 16868 1180
rect 16934 1027 16944 1180
rect 17050 1027 17060 1180
rect 17126 1027 17136 1180
rect 17242 1027 17252 1180
rect 17318 1027 17328 1180
rect 17434 1027 17444 1180
rect 17510 1027 17520 1180
rect 17626 1027 17636 1180
rect 17702 1027 17712 1180
rect 17818 1027 17828 1180
rect 17894 1027 17904 1180
rect 17940 967 18160 1214
rect 18302 1027 18312 1180
rect 18378 1027 18388 1180
rect 18494 1027 18504 1180
rect 18570 1027 18580 1180
rect 18686 1027 18696 1180
rect 18762 1027 18772 1180
rect 18878 1027 18888 1180
rect 18954 1027 18964 1180
rect 19070 1027 19080 1180
rect 19146 1027 19156 1180
rect 19262 1027 19272 1180
rect 19338 1027 19348 1180
rect 19454 1027 19464 1180
rect 19530 1027 19540 1180
rect 19646 1027 19656 1180
rect 19722 1027 19732 1180
rect 19768 967 19988 1214
rect 20130 1027 20140 1180
rect 20206 1027 20216 1180
rect 20322 1027 20332 1180
rect 20398 1027 20408 1180
rect 20514 1027 20524 1180
rect 20590 1027 20600 1180
rect 20706 1027 20716 1180
rect 20782 1027 20792 1180
rect 20898 1027 20908 1180
rect 20974 1027 20984 1180
rect 21090 1027 21100 1180
rect 21166 1027 21176 1180
rect 21282 1027 21292 1180
rect 21358 1027 21368 1180
rect 21474 1027 21484 1180
rect 21550 1027 21560 1180
rect 21596 967 21816 1214
rect 118 814 128 967
rect 194 814 204 967
rect 310 814 320 967
rect 386 814 396 967
rect 502 814 512 967
rect 578 814 588 967
rect 694 814 704 967
rect 770 814 780 967
rect 886 814 896 967
rect 962 814 972 967
rect 1078 814 1088 967
rect 1154 814 1164 967
rect 1270 814 1280 967
rect 1346 814 1356 967
rect 1462 814 1472 967
rect 1528 814 1708 967
rect 1946 814 1956 967
rect 2022 814 2032 967
rect 2138 814 2148 967
rect 2214 814 2224 967
rect 2330 814 2340 967
rect 2406 814 2416 967
rect 2522 814 2532 967
rect 2598 814 2608 967
rect 2714 814 2724 967
rect 2790 814 2800 967
rect 2906 814 2916 967
rect 2982 814 2992 967
rect 3098 814 3108 967
rect 3174 814 3184 967
rect 3290 814 3300 967
rect 3356 814 3536 967
rect 3774 814 3784 967
rect 3850 814 3860 967
rect 3966 814 3976 967
rect 4042 814 4052 967
rect 4158 814 4168 967
rect 4234 814 4244 967
rect 4350 814 4360 967
rect 4426 814 4436 967
rect 4542 814 4552 967
rect 4618 814 4628 967
rect 4734 814 4744 967
rect 4810 814 4820 967
rect 4926 814 4936 967
rect 5002 814 5012 967
rect 5118 814 5128 967
rect 5184 814 5364 967
rect 5602 814 5612 967
rect 5678 814 5688 967
rect 5794 814 5804 967
rect 5870 814 5880 967
rect 5986 814 5996 967
rect 6062 814 6072 967
rect 6178 814 6188 967
rect 6254 814 6264 967
rect 6370 814 6380 967
rect 6446 814 6456 967
rect 6562 814 6572 967
rect 6638 814 6648 967
rect 6754 814 6764 967
rect 6830 814 6840 967
rect 6946 814 6956 967
rect 7012 814 7192 967
rect 7430 814 7440 967
rect 7506 814 7516 967
rect 7622 814 7632 967
rect 7698 814 7708 967
rect 7814 814 7824 967
rect 7890 814 7900 967
rect 8006 814 8016 967
rect 8082 814 8092 967
rect 8198 814 8208 967
rect 8274 814 8284 967
rect 8390 814 8400 967
rect 8466 814 8476 967
rect 8582 814 8592 967
rect 8658 814 8668 967
rect 8774 814 8784 967
rect 8840 814 9020 967
rect 9258 814 9268 967
rect 9334 814 9344 967
rect 9450 814 9460 967
rect 9526 814 9536 967
rect 9642 814 9652 967
rect 9718 814 9728 967
rect 9834 814 9844 967
rect 9910 814 9920 967
rect 10026 814 10036 967
rect 10102 814 10112 967
rect 10218 814 10228 967
rect 10294 814 10304 967
rect 10410 814 10420 967
rect 10486 814 10496 967
rect 10602 814 10612 967
rect 10668 814 10848 967
rect 11086 814 11096 967
rect 11162 814 11172 967
rect 11278 814 11288 967
rect 11354 814 11364 967
rect 11470 814 11480 967
rect 11546 814 11556 967
rect 11662 814 11672 967
rect 11738 814 11748 967
rect 11854 814 11864 967
rect 11930 814 11940 967
rect 12046 814 12056 967
rect 12122 814 12132 967
rect 12238 814 12248 967
rect 12314 814 12324 967
rect 12430 814 12440 967
rect 12496 814 12676 967
rect 12914 814 12924 967
rect 12990 814 13000 967
rect 13106 814 13116 967
rect 13182 814 13192 967
rect 13298 814 13308 967
rect 13374 814 13384 967
rect 13490 814 13500 967
rect 13566 814 13576 967
rect 13682 814 13692 967
rect 13758 814 13768 967
rect 13874 814 13884 967
rect 13950 814 13960 967
rect 14066 814 14076 967
rect 14142 814 14152 967
rect 14258 814 14268 967
rect 14324 814 14504 967
rect 14742 814 14752 967
rect 14818 814 14828 967
rect 14934 814 14944 967
rect 15010 814 15020 967
rect 15126 814 15136 967
rect 15202 814 15212 967
rect 15318 814 15328 967
rect 15394 814 15404 967
rect 15510 814 15520 967
rect 15586 814 15596 967
rect 15702 814 15712 967
rect 15778 814 15788 967
rect 15894 814 15904 967
rect 15970 814 15980 967
rect 16086 814 16096 967
rect 16152 814 16332 967
rect 16570 814 16580 967
rect 16646 814 16656 967
rect 16762 814 16772 967
rect 16838 814 16848 967
rect 16954 814 16964 967
rect 17030 814 17040 967
rect 17146 814 17156 967
rect 17222 814 17232 967
rect 17338 814 17348 967
rect 17414 814 17424 967
rect 17530 814 17540 967
rect 17606 814 17616 967
rect 17722 814 17732 967
rect 17798 814 17808 967
rect 17914 814 17924 967
rect 17980 814 18160 967
rect 18398 814 18408 967
rect 18474 814 18484 967
rect 18590 814 18600 967
rect 18666 814 18676 967
rect 18782 814 18792 967
rect 18858 814 18868 967
rect 18974 814 18984 967
rect 19050 814 19060 967
rect 19166 814 19176 967
rect 19242 814 19252 967
rect 19358 814 19368 967
rect 19434 814 19444 967
rect 19550 814 19560 967
rect 19626 814 19636 967
rect 19742 814 19752 967
rect 19808 814 19988 967
rect 20226 814 20236 967
rect 20302 814 20312 967
rect 20418 814 20428 967
rect 20494 814 20504 967
rect 20610 814 20620 967
rect 20686 814 20696 967
rect 20802 814 20812 967
rect 20878 814 20888 967
rect 20994 814 21004 967
rect 21070 814 21080 967
rect 21186 814 21196 967
rect 21262 814 21272 967
rect 21378 814 21388 967
rect 21454 814 21464 967
rect 21570 814 21580 967
rect 21636 814 21816 967
rect 0 717 1490 776
rect 1828 717 3318 776
rect 3656 717 5146 776
rect 5484 717 6974 776
rect 7312 717 8802 776
rect 9140 717 10630 776
rect 10968 717 12458 776
rect 12796 717 14286 776
rect 14624 717 16114 776
rect 16452 717 17942 776
rect 18280 717 19770 776
rect 20108 717 21598 776
rect 0 538 1490 597
rect 1828 538 3318 597
rect 3656 538 5146 597
rect 5484 538 6974 597
rect 7312 538 8802 597
rect 9140 538 10630 597
rect 10968 538 12458 597
rect 12796 538 14286 597
rect 14624 538 16114 597
rect 16452 538 17942 597
rect 18280 538 19770 597
rect 20108 538 21598 597
rect 22 313 32 466
rect 98 313 108 466
rect 214 313 224 466
rect 290 313 300 466
rect 406 313 416 466
rect 482 313 492 466
rect 598 313 608 466
rect 674 313 684 466
rect 790 313 800 466
rect 866 313 876 466
rect 982 313 992 466
rect 1058 313 1068 466
rect 1174 313 1184 466
rect 1250 313 1260 466
rect 1366 313 1376 466
rect 1442 313 1452 466
rect 1488 253 1708 500
rect 1850 313 1860 466
rect 1926 313 1936 466
rect 2042 313 2052 466
rect 2118 313 2128 466
rect 2234 313 2244 466
rect 2310 313 2320 466
rect 2426 313 2436 466
rect 2502 313 2512 466
rect 2618 313 2628 466
rect 2694 313 2704 466
rect 2810 313 2820 466
rect 2886 313 2896 466
rect 3002 313 3012 466
rect 3078 313 3088 466
rect 3194 313 3204 466
rect 3270 313 3280 466
rect 3316 253 3536 500
rect 3678 313 3688 466
rect 3754 313 3764 466
rect 3870 313 3880 466
rect 3946 313 3956 466
rect 4062 313 4072 466
rect 4138 313 4148 466
rect 4254 313 4264 466
rect 4330 313 4340 466
rect 4446 313 4456 466
rect 4522 313 4532 466
rect 4638 313 4648 466
rect 4714 313 4724 466
rect 4830 313 4840 466
rect 4906 313 4916 466
rect 5022 313 5032 466
rect 5098 313 5108 466
rect 5144 253 5364 500
rect 5506 313 5516 466
rect 5582 313 5592 466
rect 5698 313 5708 466
rect 5774 313 5784 466
rect 5890 313 5900 466
rect 5966 313 5976 466
rect 6082 313 6092 466
rect 6158 313 6168 466
rect 6274 313 6284 466
rect 6350 313 6360 466
rect 6466 313 6476 466
rect 6542 313 6552 466
rect 6658 313 6668 466
rect 6734 313 6744 466
rect 6850 313 6860 466
rect 6926 313 6936 466
rect 6972 253 7192 500
rect 7334 313 7344 466
rect 7410 313 7420 466
rect 7526 313 7536 466
rect 7602 313 7612 466
rect 7718 313 7728 466
rect 7794 313 7804 466
rect 7910 313 7920 466
rect 7986 313 7996 466
rect 8102 313 8112 466
rect 8178 313 8188 466
rect 8294 313 8304 466
rect 8370 313 8380 466
rect 8486 313 8496 466
rect 8562 313 8572 466
rect 8678 313 8688 466
rect 8754 313 8764 466
rect 8800 253 9020 500
rect 9162 313 9172 466
rect 9238 313 9248 466
rect 9354 313 9364 466
rect 9430 313 9440 466
rect 9546 313 9556 466
rect 9622 313 9632 466
rect 9738 313 9748 466
rect 9814 313 9824 466
rect 9930 313 9940 466
rect 10006 313 10016 466
rect 10122 313 10132 466
rect 10198 313 10208 466
rect 10314 313 10324 466
rect 10390 313 10400 466
rect 10506 313 10516 466
rect 10582 313 10592 466
rect 10628 253 10848 500
rect 10990 313 11000 466
rect 11066 313 11076 466
rect 11182 313 11192 466
rect 11258 313 11268 466
rect 11374 313 11384 466
rect 11450 313 11460 466
rect 11566 313 11576 466
rect 11642 313 11652 466
rect 11758 313 11768 466
rect 11834 313 11844 466
rect 11950 313 11960 466
rect 12026 313 12036 466
rect 12142 313 12152 466
rect 12218 313 12228 466
rect 12334 313 12344 466
rect 12410 313 12420 466
rect 12456 253 12676 500
rect 12818 313 12828 466
rect 12894 313 12904 466
rect 13010 313 13020 466
rect 13086 313 13096 466
rect 13202 313 13212 466
rect 13278 313 13288 466
rect 13394 313 13404 466
rect 13470 313 13480 466
rect 13586 313 13596 466
rect 13662 313 13672 466
rect 13778 313 13788 466
rect 13854 313 13864 466
rect 13970 313 13980 466
rect 14046 313 14056 466
rect 14162 313 14172 466
rect 14238 313 14248 466
rect 14284 253 14504 500
rect 14646 313 14656 466
rect 14722 313 14732 466
rect 14838 313 14848 466
rect 14914 313 14924 466
rect 15030 313 15040 466
rect 15106 313 15116 466
rect 15222 313 15232 466
rect 15298 313 15308 466
rect 15414 313 15424 466
rect 15490 313 15500 466
rect 15606 313 15616 466
rect 15682 313 15692 466
rect 15798 313 15808 466
rect 15874 313 15884 466
rect 15990 313 16000 466
rect 16066 313 16076 466
rect 16112 253 16332 500
rect 16474 313 16484 466
rect 16550 313 16560 466
rect 16666 313 16676 466
rect 16742 313 16752 466
rect 16858 313 16868 466
rect 16934 313 16944 466
rect 17050 313 17060 466
rect 17126 313 17136 466
rect 17242 313 17252 466
rect 17318 313 17328 466
rect 17434 313 17444 466
rect 17510 313 17520 466
rect 17626 313 17636 466
rect 17702 313 17712 466
rect 17818 313 17828 466
rect 17894 313 17904 466
rect 17940 253 18160 500
rect 18302 313 18312 466
rect 18378 313 18388 466
rect 18494 313 18504 466
rect 18570 313 18580 466
rect 18686 313 18696 466
rect 18762 313 18772 466
rect 18878 313 18888 466
rect 18954 313 18964 466
rect 19070 313 19080 466
rect 19146 313 19156 466
rect 19262 313 19272 466
rect 19338 313 19348 466
rect 19454 313 19464 466
rect 19530 313 19540 466
rect 19646 313 19656 466
rect 19722 313 19732 466
rect 19768 253 19988 500
rect 20130 313 20140 466
rect 20206 313 20216 466
rect 20322 313 20332 466
rect 20398 313 20408 466
rect 20514 313 20524 466
rect 20590 313 20600 466
rect 20706 313 20716 466
rect 20782 313 20792 466
rect 20898 313 20908 466
rect 20974 313 20984 466
rect 21090 313 21100 466
rect 21166 313 21176 466
rect 21282 313 21292 466
rect 21358 313 21368 466
rect 21474 313 21484 466
rect 21550 313 21560 466
rect 21596 253 21816 500
rect 118 100 128 253
rect 194 100 204 253
rect 310 100 320 253
rect 386 100 396 253
rect 502 100 512 253
rect 578 100 588 253
rect 694 100 704 253
rect 770 100 780 253
rect 886 100 896 253
rect 962 100 972 253
rect 1078 100 1088 253
rect 1154 100 1164 253
rect 1270 100 1280 253
rect 1346 100 1356 253
rect 1462 100 1472 253
rect 1528 100 1708 253
rect 1946 100 1956 253
rect 2022 100 2032 253
rect 2138 100 2148 253
rect 2214 100 2224 253
rect 2330 100 2340 253
rect 2406 100 2416 253
rect 2522 100 2532 253
rect 2598 100 2608 253
rect 2714 100 2724 253
rect 2790 100 2800 253
rect 2906 100 2916 253
rect 2982 100 2992 253
rect 3098 100 3108 253
rect 3174 100 3184 253
rect 3290 100 3300 253
rect 3356 100 3536 253
rect 3774 100 3784 253
rect 3850 100 3860 253
rect 3966 100 3976 253
rect 4042 100 4052 253
rect 4158 100 4168 253
rect 4234 100 4244 253
rect 4350 100 4360 253
rect 4426 100 4436 253
rect 4542 100 4552 253
rect 4618 100 4628 253
rect 4734 100 4744 253
rect 4810 100 4820 253
rect 4926 100 4936 253
rect 5002 100 5012 253
rect 5118 100 5128 253
rect 5184 100 5364 253
rect 5602 100 5612 253
rect 5678 100 5688 253
rect 5794 100 5804 253
rect 5870 100 5880 253
rect 5986 100 5996 253
rect 6062 100 6072 253
rect 6178 100 6188 253
rect 6254 100 6264 253
rect 6370 100 6380 253
rect 6446 100 6456 253
rect 6562 100 6572 253
rect 6638 100 6648 253
rect 6754 100 6764 253
rect 6830 100 6840 253
rect 6946 100 6956 253
rect 7012 100 7192 253
rect 7430 100 7440 253
rect 7506 100 7516 253
rect 7622 100 7632 253
rect 7698 100 7708 253
rect 7814 100 7824 253
rect 7890 100 7900 253
rect 8006 100 8016 253
rect 8082 100 8092 253
rect 8198 100 8208 253
rect 8274 100 8284 253
rect 8390 100 8400 253
rect 8466 100 8476 253
rect 8582 100 8592 253
rect 8658 100 8668 253
rect 8774 100 8784 253
rect 8840 100 9020 253
rect 9258 100 9268 253
rect 9334 100 9344 253
rect 9450 100 9460 253
rect 9526 100 9536 253
rect 9642 100 9652 253
rect 9718 100 9728 253
rect 9834 100 9844 253
rect 9910 100 9920 253
rect 10026 100 10036 253
rect 10102 100 10112 253
rect 10218 100 10228 253
rect 10294 100 10304 253
rect 10410 100 10420 253
rect 10486 100 10496 253
rect 10602 100 10612 253
rect 10668 100 10848 253
rect 11086 100 11096 253
rect 11162 100 11172 253
rect 11278 100 11288 253
rect 11354 100 11364 253
rect 11470 100 11480 253
rect 11546 100 11556 253
rect 11662 100 11672 253
rect 11738 100 11748 253
rect 11854 100 11864 253
rect 11930 100 11940 253
rect 12046 100 12056 253
rect 12122 100 12132 253
rect 12238 100 12248 253
rect 12314 100 12324 253
rect 12430 100 12440 253
rect 12496 100 12676 253
rect 12914 100 12924 253
rect 12990 100 13000 253
rect 13106 100 13116 253
rect 13182 100 13192 253
rect 13298 100 13308 253
rect 13374 100 13384 253
rect 13490 100 13500 253
rect 13566 100 13576 253
rect 13682 100 13692 253
rect 13758 100 13768 253
rect 13874 100 13884 253
rect 13950 100 13960 253
rect 14066 100 14076 253
rect 14142 100 14152 253
rect 14258 100 14268 253
rect 14324 100 14504 253
rect 14742 100 14752 253
rect 14818 100 14828 253
rect 14934 100 14944 253
rect 15010 100 15020 253
rect 15126 100 15136 253
rect 15202 100 15212 253
rect 15318 100 15328 253
rect 15394 100 15404 253
rect 15510 100 15520 253
rect 15586 100 15596 253
rect 15702 100 15712 253
rect 15778 100 15788 253
rect 15894 100 15904 253
rect 15970 100 15980 253
rect 16086 100 16096 253
rect 16152 100 16332 253
rect 16570 100 16580 253
rect 16646 100 16656 253
rect 16762 100 16772 253
rect 16838 100 16848 253
rect 16954 100 16964 253
rect 17030 100 17040 253
rect 17146 100 17156 253
rect 17222 100 17232 253
rect 17338 100 17348 253
rect 17414 100 17424 253
rect 17530 100 17540 253
rect 17606 100 17616 253
rect 17722 100 17732 253
rect 17798 100 17808 253
rect 17914 100 17924 253
rect 17980 100 18160 253
rect 18398 100 18408 253
rect 18474 100 18484 253
rect 18590 100 18600 253
rect 18666 100 18676 253
rect 18782 100 18792 253
rect 18858 100 18868 253
rect 18974 100 18984 253
rect 19050 100 19060 253
rect 19166 100 19176 253
rect 19242 100 19252 253
rect 19358 100 19368 253
rect 19434 100 19444 253
rect 19550 100 19560 253
rect 19626 100 19636 253
rect 19742 100 19752 253
rect 19808 100 19988 253
rect 20226 100 20236 253
rect 20302 100 20312 253
rect 20418 100 20428 253
rect 20494 100 20504 253
rect 20610 100 20620 253
rect 20686 100 20696 253
rect 20802 100 20812 253
rect 20878 100 20888 253
rect 20994 100 21004 253
rect 21070 100 21080 253
rect 21186 100 21196 253
rect 21262 100 21272 253
rect 21378 100 21388 253
rect 21454 100 21464 253
rect 21570 100 21580 253
rect 21636 100 21816 253
rect 0 3 1490 62
rect 1828 3 3318 62
rect 3656 3 5146 62
rect 5484 3 6974 62
rect 7312 3 8802 62
rect 9140 3 10630 62
rect 10968 3 12458 62
rect 12796 3 14286 62
rect 14624 3 16114 62
rect 16452 3 17942 62
rect 18280 3 19770 62
rect 20108 3 21598 62
<< via1 >>
rect 32 21019 98 21172
rect 224 21019 290 21172
rect 416 21019 482 21172
rect 608 21019 674 21172
rect 800 21019 866 21172
rect 992 21019 1058 21172
rect 1184 21019 1250 21172
rect 1376 21019 1442 21172
rect 1860 21019 1926 21172
rect 2052 21019 2118 21172
rect 2244 21019 2310 21172
rect 2436 21019 2502 21172
rect 2628 21019 2694 21172
rect 2820 21019 2886 21172
rect 3012 21019 3078 21172
rect 3204 21019 3270 21172
rect 3688 21019 3754 21172
rect 3880 21019 3946 21172
rect 4072 21019 4138 21172
rect 4264 21019 4330 21172
rect 4456 21019 4522 21172
rect 4648 21019 4714 21172
rect 4840 21019 4906 21172
rect 5032 21019 5098 21172
rect 5516 21019 5582 21172
rect 5708 21019 5774 21172
rect 5900 21019 5966 21172
rect 6092 21019 6158 21172
rect 6284 21019 6350 21172
rect 6476 21019 6542 21172
rect 6668 21019 6734 21172
rect 6860 21019 6926 21172
rect 7344 21019 7410 21172
rect 7536 21019 7602 21172
rect 7728 21019 7794 21172
rect 7920 21019 7986 21172
rect 8112 21019 8178 21172
rect 8304 21019 8370 21172
rect 8496 21019 8562 21172
rect 8688 21019 8754 21172
rect 9172 21019 9238 21172
rect 9364 21019 9430 21172
rect 9556 21019 9622 21172
rect 9748 21019 9814 21172
rect 9940 21019 10006 21172
rect 10132 21019 10198 21172
rect 10324 21019 10390 21172
rect 10516 21019 10582 21172
rect 11000 21019 11066 21172
rect 11192 21019 11258 21172
rect 11384 21019 11450 21172
rect 11576 21019 11642 21172
rect 11768 21019 11834 21172
rect 11960 21019 12026 21172
rect 12152 21019 12218 21172
rect 12344 21019 12410 21172
rect 12828 21019 12894 21172
rect 13020 21019 13086 21172
rect 13212 21019 13278 21172
rect 13404 21019 13470 21172
rect 13596 21019 13662 21172
rect 13788 21019 13854 21172
rect 13980 21019 14046 21172
rect 14172 21019 14238 21172
rect 14656 21019 14722 21172
rect 14848 21019 14914 21172
rect 15040 21019 15106 21172
rect 15232 21019 15298 21172
rect 15424 21019 15490 21172
rect 15616 21019 15682 21172
rect 15808 21019 15874 21172
rect 16000 21019 16066 21172
rect 16484 21019 16550 21172
rect 16676 21019 16742 21172
rect 16868 21019 16934 21172
rect 17060 21019 17126 21172
rect 17252 21019 17318 21172
rect 17444 21019 17510 21172
rect 17636 21019 17702 21172
rect 17828 21019 17894 21172
rect 18312 21019 18378 21172
rect 18504 21019 18570 21172
rect 18696 21019 18762 21172
rect 18888 21019 18954 21172
rect 19080 21019 19146 21172
rect 19272 21019 19338 21172
rect 19464 21019 19530 21172
rect 19656 21019 19722 21172
rect 20140 21019 20206 21172
rect 20332 21019 20398 21172
rect 20524 21019 20590 21172
rect 20716 21019 20782 21172
rect 20908 21019 20974 21172
rect 21100 21019 21166 21172
rect 21292 21019 21358 21172
rect 21484 21019 21550 21172
rect 128 20806 194 20959
rect 320 20806 386 20959
rect 512 20806 578 20959
rect 704 20806 770 20959
rect 896 20806 962 20959
rect 1088 20806 1154 20959
rect 1280 20806 1346 20959
rect 1472 20806 1528 20959
rect 1956 20806 2022 20959
rect 2148 20806 2214 20959
rect 2340 20806 2406 20959
rect 2532 20806 2598 20959
rect 2724 20806 2790 20959
rect 2916 20806 2982 20959
rect 3108 20806 3174 20959
rect 3300 20806 3356 20959
rect 3784 20806 3850 20959
rect 3976 20806 4042 20959
rect 4168 20806 4234 20959
rect 4360 20806 4426 20959
rect 4552 20806 4618 20959
rect 4744 20806 4810 20959
rect 4936 20806 5002 20959
rect 5128 20806 5184 20959
rect 5612 20806 5678 20959
rect 5804 20806 5870 20959
rect 5996 20806 6062 20959
rect 6188 20806 6254 20959
rect 6380 20806 6446 20959
rect 6572 20806 6638 20959
rect 6764 20806 6830 20959
rect 6956 20806 7012 20959
rect 7440 20806 7506 20959
rect 7632 20806 7698 20959
rect 7824 20806 7890 20959
rect 8016 20806 8082 20959
rect 8208 20806 8274 20959
rect 8400 20806 8466 20959
rect 8592 20806 8658 20959
rect 8784 20806 8840 20959
rect 9268 20806 9334 20959
rect 9460 20806 9526 20959
rect 9652 20806 9718 20959
rect 9844 20806 9910 20959
rect 10036 20806 10102 20959
rect 10228 20806 10294 20959
rect 10420 20806 10486 20959
rect 10612 20806 10668 20959
rect 11096 20806 11162 20959
rect 11288 20806 11354 20959
rect 11480 20806 11546 20959
rect 11672 20806 11738 20959
rect 11864 20806 11930 20959
rect 12056 20806 12122 20959
rect 12248 20806 12314 20959
rect 12440 20806 12496 20959
rect 12924 20806 12990 20959
rect 13116 20806 13182 20959
rect 13308 20806 13374 20959
rect 13500 20806 13566 20959
rect 13692 20806 13758 20959
rect 13884 20806 13950 20959
rect 14076 20806 14142 20959
rect 14268 20806 14324 20959
rect 14752 20806 14818 20959
rect 14944 20806 15010 20959
rect 15136 20806 15202 20959
rect 15328 20806 15394 20959
rect 15520 20806 15586 20959
rect 15712 20806 15778 20959
rect 15904 20806 15970 20959
rect 16096 20806 16152 20959
rect 16580 20806 16646 20959
rect 16772 20806 16838 20959
rect 16964 20806 17030 20959
rect 17156 20806 17222 20959
rect 17348 20806 17414 20959
rect 17540 20806 17606 20959
rect 17732 20806 17798 20959
rect 17924 20806 17980 20959
rect 18408 20806 18474 20959
rect 18600 20806 18666 20959
rect 18792 20806 18858 20959
rect 18984 20806 19050 20959
rect 19176 20806 19242 20959
rect 19368 20806 19434 20959
rect 19560 20806 19626 20959
rect 19752 20806 19808 20959
rect 20236 20806 20302 20959
rect 20428 20806 20494 20959
rect 20620 20806 20686 20959
rect 20812 20806 20878 20959
rect 21004 20806 21070 20959
rect 21196 20806 21262 20959
rect 21388 20806 21454 20959
rect 21580 20806 21636 20959
rect 32 20305 98 20458
rect 224 20305 290 20458
rect 416 20305 482 20458
rect 608 20305 674 20458
rect 800 20305 866 20458
rect 992 20305 1058 20458
rect 1184 20305 1250 20458
rect 1376 20305 1442 20458
rect 1860 20305 1926 20458
rect 2052 20305 2118 20458
rect 2244 20305 2310 20458
rect 2436 20305 2502 20458
rect 2628 20305 2694 20458
rect 2820 20305 2886 20458
rect 3012 20305 3078 20458
rect 3204 20305 3270 20458
rect 3688 20305 3754 20458
rect 3880 20305 3946 20458
rect 4072 20305 4138 20458
rect 4264 20305 4330 20458
rect 4456 20305 4522 20458
rect 4648 20305 4714 20458
rect 4840 20305 4906 20458
rect 5032 20305 5098 20458
rect 5516 20305 5582 20458
rect 5708 20305 5774 20458
rect 5900 20305 5966 20458
rect 6092 20305 6158 20458
rect 6284 20305 6350 20458
rect 6476 20305 6542 20458
rect 6668 20305 6734 20458
rect 6860 20305 6926 20458
rect 7344 20305 7410 20458
rect 7536 20305 7602 20458
rect 7728 20305 7794 20458
rect 7920 20305 7986 20458
rect 8112 20305 8178 20458
rect 8304 20305 8370 20458
rect 8496 20305 8562 20458
rect 8688 20305 8754 20458
rect 9172 20305 9238 20458
rect 9364 20305 9430 20458
rect 9556 20305 9622 20458
rect 9748 20305 9814 20458
rect 9940 20305 10006 20458
rect 10132 20305 10198 20458
rect 10324 20305 10390 20458
rect 10516 20305 10582 20458
rect 11000 20305 11066 20458
rect 11192 20305 11258 20458
rect 11384 20305 11450 20458
rect 11576 20305 11642 20458
rect 11768 20305 11834 20458
rect 11960 20305 12026 20458
rect 12152 20305 12218 20458
rect 12344 20305 12410 20458
rect 12828 20305 12894 20458
rect 13020 20305 13086 20458
rect 13212 20305 13278 20458
rect 13404 20305 13470 20458
rect 13596 20305 13662 20458
rect 13788 20305 13854 20458
rect 13980 20305 14046 20458
rect 14172 20305 14238 20458
rect 14656 20305 14722 20458
rect 14848 20305 14914 20458
rect 15040 20305 15106 20458
rect 15232 20305 15298 20458
rect 15424 20305 15490 20458
rect 15616 20305 15682 20458
rect 15808 20305 15874 20458
rect 16000 20305 16066 20458
rect 16484 20305 16550 20458
rect 16676 20305 16742 20458
rect 16868 20305 16934 20458
rect 17060 20305 17126 20458
rect 17252 20305 17318 20458
rect 17444 20305 17510 20458
rect 17636 20305 17702 20458
rect 17828 20305 17894 20458
rect 18312 20305 18378 20458
rect 18504 20305 18570 20458
rect 18696 20305 18762 20458
rect 18888 20305 18954 20458
rect 19080 20305 19146 20458
rect 19272 20305 19338 20458
rect 19464 20305 19530 20458
rect 19656 20305 19722 20458
rect 20140 20305 20206 20458
rect 20332 20305 20398 20458
rect 20524 20305 20590 20458
rect 20716 20305 20782 20458
rect 20908 20305 20974 20458
rect 21100 20305 21166 20458
rect 21292 20305 21358 20458
rect 21484 20305 21550 20458
rect 128 20092 194 20245
rect 320 20092 386 20245
rect 512 20092 578 20245
rect 704 20092 770 20245
rect 896 20092 962 20245
rect 1088 20092 1154 20245
rect 1280 20092 1346 20245
rect 1472 20092 1528 20245
rect 1956 20092 2022 20245
rect 2148 20092 2214 20245
rect 2340 20092 2406 20245
rect 2532 20092 2598 20245
rect 2724 20092 2790 20245
rect 2916 20092 2982 20245
rect 3108 20092 3174 20245
rect 3300 20092 3356 20245
rect 3784 20092 3850 20245
rect 3976 20092 4042 20245
rect 4168 20092 4234 20245
rect 4360 20092 4426 20245
rect 4552 20092 4618 20245
rect 4744 20092 4810 20245
rect 4936 20092 5002 20245
rect 5128 20092 5184 20245
rect 5612 20092 5678 20245
rect 5804 20092 5870 20245
rect 5996 20092 6062 20245
rect 6188 20092 6254 20245
rect 6380 20092 6446 20245
rect 6572 20092 6638 20245
rect 6764 20092 6830 20245
rect 6956 20092 7012 20245
rect 7440 20092 7506 20245
rect 7632 20092 7698 20245
rect 7824 20092 7890 20245
rect 8016 20092 8082 20245
rect 8208 20092 8274 20245
rect 8400 20092 8466 20245
rect 8592 20092 8658 20245
rect 8784 20092 8840 20245
rect 9268 20092 9334 20245
rect 9460 20092 9526 20245
rect 9652 20092 9718 20245
rect 9844 20092 9910 20245
rect 10036 20092 10102 20245
rect 10228 20092 10294 20245
rect 10420 20092 10486 20245
rect 10612 20092 10668 20245
rect 11096 20092 11162 20245
rect 11288 20092 11354 20245
rect 11480 20092 11546 20245
rect 11672 20092 11738 20245
rect 11864 20092 11930 20245
rect 12056 20092 12122 20245
rect 12248 20092 12314 20245
rect 12440 20092 12496 20245
rect 12924 20092 12990 20245
rect 13116 20092 13182 20245
rect 13308 20092 13374 20245
rect 13500 20092 13566 20245
rect 13692 20092 13758 20245
rect 13884 20092 13950 20245
rect 14076 20092 14142 20245
rect 14268 20092 14324 20245
rect 14752 20092 14818 20245
rect 14944 20092 15010 20245
rect 15136 20092 15202 20245
rect 15328 20092 15394 20245
rect 15520 20092 15586 20245
rect 15712 20092 15778 20245
rect 15904 20092 15970 20245
rect 16096 20092 16152 20245
rect 16580 20092 16646 20245
rect 16772 20092 16838 20245
rect 16964 20092 17030 20245
rect 17156 20092 17222 20245
rect 17348 20092 17414 20245
rect 17540 20092 17606 20245
rect 17732 20092 17798 20245
rect 17924 20092 17980 20245
rect 18408 20092 18474 20245
rect 18600 20092 18666 20245
rect 18792 20092 18858 20245
rect 18984 20092 19050 20245
rect 19176 20092 19242 20245
rect 19368 20092 19434 20245
rect 19560 20092 19626 20245
rect 19752 20092 19808 20245
rect 20236 20092 20302 20245
rect 20428 20092 20494 20245
rect 20620 20092 20686 20245
rect 20812 20092 20878 20245
rect 21004 20092 21070 20245
rect 21196 20092 21262 20245
rect 21388 20092 21454 20245
rect 21580 20092 21636 20245
rect 32 19591 98 19744
rect 224 19591 290 19744
rect 416 19591 482 19744
rect 608 19591 674 19744
rect 800 19591 866 19744
rect 992 19591 1058 19744
rect 1184 19591 1250 19744
rect 1376 19591 1442 19744
rect 1860 19591 1926 19744
rect 2052 19591 2118 19744
rect 2244 19591 2310 19744
rect 2436 19591 2502 19744
rect 2628 19591 2694 19744
rect 2820 19591 2886 19744
rect 3012 19591 3078 19744
rect 3204 19591 3270 19744
rect 3688 19591 3754 19744
rect 3880 19591 3946 19744
rect 4072 19591 4138 19744
rect 4264 19591 4330 19744
rect 4456 19591 4522 19744
rect 4648 19591 4714 19744
rect 4840 19591 4906 19744
rect 5032 19591 5098 19744
rect 5516 19591 5582 19744
rect 5708 19591 5774 19744
rect 5900 19591 5966 19744
rect 6092 19591 6158 19744
rect 6284 19591 6350 19744
rect 6476 19591 6542 19744
rect 6668 19591 6734 19744
rect 6860 19591 6926 19744
rect 7344 19591 7410 19744
rect 7536 19591 7602 19744
rect 7728 19591 7794 19744
rect 7920 19591 7986 19744
rect 8112 19591 8178 19744
rect 8304 19591 8370 19744
rect 8496 19591 8562 19744
rect 8688 19591 8754 19744
rect 9172 19591 9238 19744
rect 9364 19591 9430 19744
rect 9556 19591 9622 19744
rect 9748 19591 9814 19744
rect 9940 19591 10006 19744
rect 10132 19591 10198 19744
rect 10324 19591 10390 19744
rect 10516 19591 10582 19744
rect 11000 19591 11066 19744
rect 11192 19591 11258 19744
rect 11384 19591 11450 19744
rect 11576 19591 11642 19744
rect 11768 19591 11834 19744
rect 11960 19591 12026 19744
rect 12152 19591 12218 19744
rect 12344 19591 12410 19744
rect 12828 19591 12894 19744
rect 13020 19591 13086 19744
rect 13212 19591 13278 19744
rect 13404 19591 13470 19744
rect 13596 19591 13662 19744
rect 13788 19591 13854 19744
rect 13980 19591 14046 19744
rect 14172 19591 14238 19744
rect 14656 19591 14722 19744
rect 14848 19591 14914 19744
rect 15040 19591 15106 19744
rect 15232 19591 15298 19744
rect 15424 19591 15490 19744
rect 15616 19591 15682 19744
rect 15808 19591 15874 19744
rect 16000 19591 16066 19744
rect 16484 19591 16550 19744
rect 16676 19591 16742 19744
rect 16868 19591 16934 19744
rect 17060 19591 17126 19744
rect 17252 19591 17318 19744
rect 17444 19591 17510 19744
rect 17636 19591 17702 19744
rect 17828 19591 17894 19744
rect 18312 19591 18378 19744
rect 18504 19591 18570 19744
rect 18696 19591 18762 19744
rect 18888 19591 18954 19744
rect 19080 19591 19146 19744
rect 19272 19591 19338 19744
rect 19464 19591 19530 19744
rect 19656 19591 19722 19744
rect 20140 19591 20206 19744
rect 20332 19591 20398 19744
rect 20524 19591 20590 19744
rect 20716 19591 20782 19744
rect 20908 19591 20974 19744
rect 21100 19591 21166 19744
rect 21292 19591 21358 19744
rect 21484 19591 21550 19744
rect 128 19378 194 19531
rect 320 19378 386 19531
rect 512 19378 578 19531
rect 704 19378 770 19531
rect 896 19378 962 19531
rect 1088 19378 1154 19531
rect 1280 19378 1346 19531
rect 1472 19378 1528 19531
rect 1956 19378 2022 19531
rect 2148 19378 2214 19531
rect 2340 19378 2406 19531
rect 2532 19378 2598 19531
rect 2724 19378 2790 19531
rect 2916 19378 2982 19531
rect 3108 19378 3174 19531
rect 3300 19378 3356 19531
rect 3784 19378 3850 19531
rect 3976 19378 4042 19531
rect 4168 19378 4234 19531
rect 4360 19378 4426 19531
rect 4552 19378 4618 19531
rect 4744 19378 4810 19531
rect 4936 19378 5002 19531
rect 5128 19378 5184 19531
rect 5612 19378 5678 19531
rect 5804 19378 5870 19531
rect 5996 19378 6062 19531
rect 6188 19378 6254 19531
rect 6380 19378 6446 19531
rect 6572 19378 6638 19531
rect 6764 19378 6830 19531
rect 6956 19378 7012 19531
rect 7440 19378 7506 19531
rect 7632 19378 7698 19531
rect 7824 19378 7890 19531
rect 8016 19378 8082 19531
rect 8208 19378 8274 19531
rect 8400 19378 8466 19531
rect 8592 19378 8658 19531
rect 8784 19378 8840 19531
rect 9268 19378 9334 19531
rect 9460 19378 9526 19531
rect 9652 19378 9718 19531
rect 9844 19378 9910 19531
rect 10036 19378 10102 19531
rect 10228 19378 10294 19531
rect 10420 19378 10486 19531
rect 10612 19378 10668 19531
rect 11096 19378 11162 19531
rect 11288 19378 11354 19531
rect 11480 19378 11546 19531
rect 11672 19378 11738 19531
rect 11864 19378 11930 19531
rect 12056 19378 12122 19531
rect 12248 19378 12314 19531
rect 12440 19378 12496 19531
rect 12924 19378 12990 19531
rect 13116 19378 13182 19531
rect 13308 19378 13374 19531
rect 13500 19378 13566 19531
rect 13692 19378 13758 19531
rect 13884 19378 13950 19531
rect 14076 19378 14142 19531
rect 14268 19378 14324 19531
rect 14752 19378 14818 19531
rect 14944 19378 15010 19531
rect 15136 19378 15202 19531
rect 15328 19378 15394 19531
rect 15520 19378 15586 19531
rect 15712 19378 15778 19531
rect 15904 19378 15970 19531
rect 16096 19378 16152 19531
rect 16580 19378 16646 19531
rect 16772 19378 16838 19531
rect 16964 19378 17030 19531
rect 17156 19378 17222 19531
rect 17348 19378 17414 19531
rect 17540 19378 17606 19531
rect 17732 19378 17798 19531
rect 17924 19378 17980 19531
rect 18408 19378 18474 19531
rect 18600 19378 18666 19531
rect 18792 19378 18858 19531
rect 18984 19378 19050 19531
rect 19176 19378 19242 19531
rect 19368 19378 19434 19531
rect 19560 19378 19626 19531
rect 19752 19378 19808 19531
rect 20236 19378 20302 19531
rect 20428 19378 20494 19531
rect 20620 19378 20686 19531
rect 20812 19378 20878 19531
rect 21004 19378 21070 19531
rect 21196 19378 21262 19531
rect 21388 19378 21454 19531
rect 21580 19378 21636 19531
rect 32 18877 98 19030
rect 224 18877 290 19030
rect 416 18877 482 19030
rect 608 18877 674 19030
rect 800 18877 866 19030
rect 992 18877 1058 19030
rect 1184 18877 1250 19030
rect 1376 18877 1442 19030
rect 1860 18877 1926 19030
rect 2052 18877 2118 19030
rect 2244 18877 2310 19030
rect 2436 18877 2502 19030
rect 2628 18877 2694 19030
rect 2820 18877 2886 19030
rect 3012 18877 3078 19030
rect 3204 18877 3270 19030
rect 3688 18877 3754 19030
rect 3880 18877 3946 19030
rect 4072 18877 4138 19030
rect 4264 18877 4330 19030
rect 4456 18877 4522 19030
rect 4648 18877 4714 19030
rect 4840 18877 4906 19030
rect 5032 18877 5098 19030
rect 5516 18877 5582 19030
rect 5708 18877 5774 19030
rect 5900 18877 5966 19030
rect 6092 18877 6158 19030
rect 6284 18877 6350 19030
rect 6476 18877 6542 19030
rect 6668 18877 6734 19030
rect 6860 18877 6926 19030
rect 7344 18877 7410 19030
rect 7536 18877 7602 19030
rect 7728 18877 7794 19030
rect 7920 18877 7986 19030
rect 8112 18877 8178 19030
rect 8304 18877 8370 19030
rect 8496 18877 8562 19030
rect 8688 18877 8754 19030
rect 9172 18877 9238 19030
rect 9364 18877 9430 19030
rect 9556 18877 9622 19030
rect 9748 18877 9814 19030
rect 9940 18877 10006 19030
rect 10132 18877 10198 19030
rect 10324 18877 10390 19030
rect 10516 18877 10582 19030
rect 11000 18877 11066 19030
rect 11192 18877 11258 19030
rect 11384 18877 11450 19030
rect 11576 18877 11642 19030
rect 11768 18877 11834 19030
rect 11960 18877 12026 19030
rect 12152 18877 12218 19030
rect 12344 18877 12410 19030
rect 12828 18877 12894 19030
rect 13020 18877 13086 19030
rect 13212 18877 13278 19030
rect 13404 18877 13470 19030
rect 13596 18877 13662 19030
rect 13788 18877 13854 19030
rect 13980 18877 14046 19030
rect 14172 18877 14238 19030
rect 14656 18877 14722 19030
rect 14848 18877 14914 19030
rect 15040 18877 15106 19030
rect 15232 18877 15298 19030
rect 15424 18877 15490 19030
rect 15616 18877 15682 19030
rect 15808 18877 15874 19030
rect 16000 18877 16066 19030
rect 16484 18877 16550 19030
rect 16676 18877 16742 19030
rect 16868 18877 16934 19030
rect 17060 18877 17126 19030
rect 17252 18877 17318 19030
rect 17444 18877 17510 19030
rect 17636 18877 17702 19030
rect 17828 18877 17894 19030
rect 18312 18877 18378 19030
rect 18504 18877 18570 19030
rect 18696 18877 18762 19030
rect 18888 18877 18954 19030
rect 19080 18877 19146 19030
rect 19272 18877 19338 19030
rect 19464 18877 19530 19030
rect 19656 18877 19722 19030
rect 20140 18877 20206 19030
rect 20332 18877 20398 19030
rect 20524 18877 20590 19030
rect 20716 18877 20782 19030
rect 20908 18877 20974 19030
rect 21100 18877 21166 19030
rect 21292 18877 21358 19030
rect 21484 18877 21550 19030
rect 128 18664 194 18817
rect 320 18664 386 18817
rect 512 18664 578 18817
rect 704 18664 770 18817
rect 896 18664 962 18817
rect 1088 18664 1154 18817
rect 1280 18664 1346 18817
rect 1472 18664 1528 18817
rect 1956 18664 2022 18817
rect 2148 18664 2214 18817
rect 2340 18664 2406 18817
rect 2532 18664 2598 18817
rect 2724 18664 2790 18817
rect 2916 18664 2982 18817
rect 3108 18664 3174 18817
rect 3300 18664 3356 18817
rect 3784 18664 3850 18817
rect 3976 18664 4042 18817
rect 4168 18664 4234 18817
rect 4360 18664 4426 18817
rect 4552 18664 4618 18817
rect 4744 18664 4810 18817
rect 4936 18664 5002 18817
rect 5128 18664 5184 18817
rect 5612 18664 5678 18817
rect 5804 18664 5870 18817
rect 5996 18664 6062 18817
rect 6188 18664 6254 18817
rect 6380 18664 6446 18817
rect 6572 18664 6638 18817
rect 6764 18664 6830 18817
rect 6956 18664 7012 18817
rect 7440 18664 7506 18817
rect 7632 18664 7698 18817
rect 7824 18664 7890 18817
rect 8016 18664 8082 18817
rect 8208 18664 8274 18817
rect 8400 18664 8466 18817
rect 8592 18664 8658 18817
rect 8784 18664 8840 18817
rect 9268 18664 9334 18817
rect 9460 18664 9526 18817
rect 9652 18664 9718 18817
rect 9844 18664 9910 18817
rect 10036 18664 10102 18817
rect 10228 18664 10294 18817
rect 10420 18664 10486 18817
rect 10612 18664 10668 18817
rect 11096 18664 11162 18817
rect 11288 18664 11354 18817
rect 11480 18664 11546 18817
rect 11672 18664 11738 18817
rect 11864 18664 11930 18817
rect 12056 18664 12122 18817
rect 12248 18664 12314 18817
rect 12440 18664 12496 18817
rect 12924 18664 12990 18817
rect 13116 18664 13182 18817
rect 13308 18664 13374 18817
rect 13500 18664 13566 18817
rect 13692 18664 13758 18817
rect 13884 18664 13950 18817
rect 14076 18664 14142 18817
rect 14268 18664 14324 18817
rect 14752 18664 14818 18817
rect 14944 18664 15010 18817
rect 15136 18664 15202 18817
rect 15328 18664 15394 18817
rect 15520 18664 15586 18817
rect 15712 18664 15778 18817
rect 15904 18664 15970 18817
rect 16096 18664 16152 18817
rect 16580 18664 16646 18817
rect 16772 18664 16838 18817
rect 16964 18664 17030 18817
rect 17156 18664 17222 18817
rect 17348 18664 17414 18817
rect 17540 18664 17606 18817
rect 17732 18664 17798 18817
rect 17924 18664 17980 18817
rect 18408 18664 18474 18817
rect 18600 18664 18666 18817
rect 18792 18664 18858 18817
rect 18984 18664 19050 18817
rect 19176 18664 19242 18817
rect 19368 18664 19434 18817
rect 19560 18664 19626 18817
rect 19752 18664 19808 18817
rect 20236 18664 20302 18817
rect 20428 18664 20494 18817
rect 20620 18664 20686 18817
rect 20812 18664 20878 18817
rect 21004 18664 21070 18817
rect 21196 18664 21262 18817
rect 21388 18664 21454 18817
rect 21580 18664 21636 18817
rect 32 18163 98 18316
rect 224 18163 290 18316
rect 416 18163 482 18316
rect 608 18163 674 18316
rect 800 18163 866 18316
rect 992 18163 1058 18316
rect 1184 18163 1250 18316
rect 1376 18163 1442 18316
rect 1860 18163 1926 18316
rect 2052 18163 2118 18316
rect 2244 18163 2310 18316
rect 2436 18163 2502 18316
rect 2628 18163 2694 18316
rect 2820 18163 2886 18316
rect 3012 18163 3078 18316
rect 3204 18163 3270 18316
rect 3688 18163 3754 18316
rect 3880 18163 3946 18316
rect 4072 18163 4138 18316
rect 4264 18163 4330 18316
rect 4456 18163 4522 18316
rect 4648 18163 4714 18316
rect 4840 18163 4906 18316
rect 5032 18163 5098 18316
rect 5516 18163 5582 18316
rect 5708 18163 5774 18316
rect 5900 18163 5966 18316
rect 6092 18163 6158 18316
rect 6284 18163 6350 18316
rect 6476 18163 6542 18316
rect 6668 18163 6734 18316
rect 6860 18163 6926 18316
rect 7344 18163 7410 18316
rect 7536 18163 7602 18316
rect 7728 18163 7794 18316
rect 7920 18163 7986 18316
rect 8112 18163 8178 18316
rect 8304 18163 8370 18316
rect 8496 18163 8562 18316
rect 8688 18163 8754 18316
rect 9172 18163 9238 18316
rect 9364 18163 9430 18316
rect 9556 18163 9622 18316
rect 9748 18163 9814 18316
rect 9940 18163 10006 18316
rect 10132 18163 10198 18316
rect 10324 18163 10390 18316
rect 10516 18163 10582 18316
rect 11000 18163 11066 18316
rect 11192 18163 11258 18316
rect 11384 18163 11450 18316
rect 11576 18163 11642 18316
rect 11768 18163 11834 18316
rect 11960 18163 12026 18316
rect 12152 18163 12218 18316
rect 12344 18163 12410 18316
rect 12828 18163 12894 18316
rect 13020 18163 13086 18316
rect 13212 18163 13278 18316
rect 13404 18163 13470 18316
rect 13596 18163 13662 18316
rect 13788 18163 13854 18316
rect 13980 18163 14046 18316
rect 14172 18163 14238 18316
rect 14656 18163 14722 18316
rect 14848 18163 14914 18316
rect 15040 18163 15106 18316
rect 15232 18163 15298 18316
rect 15424 18163 15490 18316
rect 15616 18163 15682 18316
rect 15808 18163 15874 18316
rect 16000 18163 16066 18316
rect 16484 18163 16550 18316
rect 16676 18163 16742 18316
rect 16868 18163 16934 18316
rect 17060 18163 17126 18316
rect 17252 18163 17318 18316
rect 17444 18163 17510 18316
rect 17636 18163 17702 18316
rect 17828 18163 17894 18316
rect 18312 18163 18378 18316
rect 18504 18163 18570 18316
rect 18696 18163 18762 18316
rect 18888 18163 18954 18316
rect 19080 18163 19146 18316
rect 19272 18163 19338 18316
rect 19464 18163 19530 18316
rect 19656 18163 19722 18316
rect 20140 18163 20206 18316
rect 20332 18163 20398 18316
rect 20524 18163 20590 18316
rect 20716 18163 20782 18316
rect 20908 18163 20974 18316
rect 21100 18163 21166 18316
rect 21292 18163 21358 18316
rect 21484 18163 21550 18316
rect 128 17950 194 18103
rect 320 17950 386 18103
rect 512 17950 578 18103
rect 704 17950 770 18103
rect 896 17950 962 18103
rect 1088 17950 1154 18103
rect 1280 17950 1346 18103
rect 1472 17950 1528 18103
rect 1956 17950 2022 18103
rect 2148 17950 2214 18103
rect 2340 17950 2406 18103
rect 2532 17950 2598 18103
rect 2724 17950 2790 18103
rect 2916 17950 2982 18103
rect 3108 17950 3174 18103
rect 3300 17950 3356 18103
rect 3784 17950 3850 18103
rect 3976 17950 4042 18103
rect 4168 17950 4234 18103
rect 4360 17950 4426 18103
rect 4552 17950 4618 18103
rect 4744 17950 4810 18103
rect 4936 17950 5002 18103
rect 5128 17950 5184 18103
rect 5612 17950 5678 18103
rect 5804 17950 5870 18103
rect 5996 17950 6062 18103
rect 6188 17950 6254 18103
rect 6380 17950 6446 18103
rect 6572 17950 6638 18103
rect 6764 17950 6830 18103
rect 6956 17950 7012 18103
rect 7440 17950 7506 18103
rect 7632 17950 7698 18103
rect 7824 17950 7890 18103
rect 8016 17950 8082 18103
rect 8208 17950 8274 18103
rect 8400 17950 8466 18103
rect 8592 17950 8658 18103
rect 8784 17950 8840 18103
rect 9268 17950 9334 18103
rect 9460 17950 9526 18103
rect 9652 17950 9718 18103
rect 9844 17950 9910 18103
rect 10036 17950 10102 18103
rect 10228 17950 10294 18103
rect 10420 17950 10486 18103
rect 10612 17950 10668 18103
rect 11096 17950 11162 18103
rect 11288 17950 11354 18103
rect 11480 17950 11546 18103
rect 11672 17950 11738 18103
rect 11864 17950 11930 18103
rect 12056 17950 12122 18103
rect 12248 17950 12314 18103
rect 12440 17950 12496 18103
rect 12924 17950 12990 18103
rect 13116 17950 13182 18103
rect 13308 17950 13374 18103
rect 13500 17950 13566 18103
rect 13692 17950 13758 18103
rect 13884 17950 13950 18103
rect 14076 17950 14142 18103
rect 14268 17950 14324 18103
rect 14752 17950 14818 18103
rect 14944 17950 15010 18103
rect 15136 17950 15202 18103
rect 15328 17950 15394 18103
rect 15520 17950 15586 18103
rect 15712 17950 15778 18103
rect 15904 17950 15970 18103
rect 16096 17950 16152 18103
rect 16580 17950 16646 18103
rect 16772 17950 16838 18103
rect 16964 17950 17030 18103
rect 17156 17950 17222 18103
rect 17348 17950 17414 18103
rect 17540 17950 17606 18103
rect 17732 17950 17798 18103
rect 17924 17950 17980 18103
rect 18408 17950 18474 18103
rect 18600 17950 18666 18103
rect 18792 17950 18858 18103
rect 18984 17950 19050 18103
rect 19176 17950 19242 18103
rect 19368 17950 19434 18103
rect 19560 17950 19626 18103
rect 19752 17950 19808 18103
rect 20236 17950 20302 18103
rect 20428 17950 20494 18103
rect 20620 17950 20686 18103
rect 20812 17950 20878 18103
rect 21004 17950 21070 18103
rect 21196 17950 21262 18103
rect 21388 17950 21454 18103
rect 21580 17950 21636 18103
rect 32 17449 98 17602
rect 224 17449 290 17602
rect 416 17449 482 17602
rect 608 17449 674 17602
rect 800 17449 866 17602
rect 992 17449 1058 17602
rect 1184 17449 1250 17602
rect 1376 17449 1442 17602
rect 1860 17449 1926 17602
rect 2052 17449 2118 17602
rect 2244 17449 2310 17602
rect 2436 17449 2502 17602
rect 2628 17449 2694 17602
rect 2820 17449 2886 17602
rect 3012 17449 3078 17602
rect 3204 17449 3270 17602
rect 3688 17449 3754 17602
rect 3880 17449 3946 17602
rect 4072 17449 4138 17602
rect 4264 17449 4330 17602
rect 4456 17449 4522 17602
rect 4648 17449 4714 17602
rect 4840 17449 4906 17602
rect 5032 17449 5098 17602
rect 5516 17449 5582 17602
rect 5708 17449 5774 17602
rect 5900 17449 5966 17602
rect 6092 17449 6158 17602
rect 6284 17449 6350 17602
rect 6476 17449 6542 17602
rect 6668 17449 6734 17602
rect 6860 17449 6926 17602
rect 7344 17449 7410 17602
rect 7536 17449 7602 17602
rect 7728 17449 7794 17602
rect 7920 17449 7986 17602
rect 8112 17449 8178 17602
rect 8304 17449 8370 17602
rect 8496 17449 8562 17602
rect 8688 17449 8754 17602
rect 9172 17449 9238 17602
rect 9364 17449 9430 17602
rect 9556 17449 9622 17602
rect 9748 17449 9814 17602
rect 9940 17449 10006 17602
rect 10132 17449 10198 17602
rect 10324 17449 10390 17602
rect 10516 17449 10582 17602
rect 11000 17449 11066 17602
rect 11192 17449 11258 17602
rect 11384 17449 11450 17602
rect 11576 17449 11642 17602
rect 11768 17449 11834 17602
rect 11960 17449 12026 17602
rect 12152 17449 12218 17602
rect 12344 17449 12410 17602
rect 12828 17449 12894 17602
rect 13020 17449 13086 17602
rect 13212 17449 13278 17602
rect 13404 17449 13470 17602
rect 13596 17449 13662 17602
rect 13788 17449 13854 17602
rect 13980 17449 14046 17602
rect 14172 17449 14238 17602
rect 14656 17449 14722 17602
rect 14848 17449 14914 17602
rect 15040 17449 15106 17602
rect 15232 17449 15298 17602
rect 15424 17449 15490 17602
rect 15616 17449 15682 17602
rect 15808 17449 15874 17602
rect 16000 17449 16066 17602
rect 16484 17449 16550 17602
rect 16676 17449 16742 17602
rect 16868 17449 16934 17602
rect 17060 17449 17126 17602
rect 17252 17449 17318 17602
rect 17444 17449 17510 17602
rect 17636 17449 17702 17602
rect 17828 17449 17894 17602
rect 18312 17449 18378 17602
rect 18504 17449 18570 17602
rect 18696 17449 18762 17602
rect 18888 17449 18954 17602
rect 19080 17449 19146 17602
rect 19272 17449 19338 17602
rect 19464 17449 19530 17602
rect 19656 17449 19722 17602
rect 20140 17449 20206 17602
rect 20332 17449 20398 17602
rect 20524 17449 20590 17602
rect 20716 17449 20782 17602
rect 20908 17449 20974 17602
rect 21100 17449 21166 17602
rect 21292 17449 21358 17602
rect 21484 17449 21550 17602
rect 128 17236 194 17389
rect 320 17236 386 17389
rect 512 17236 578 17389
rect 704 17236 770 17389
rect 896 17236 962 17389
rect 1088 17236 1154 17389
rect 1280 17236 1346 17389
rect 1472 17236 1528 17389
rect 1956 17236 2022 17389
rect 2148 17236 2214 17389
rect 2340 17236 2406 17389
rect 2532 17236 2598 17389
rect 2724 17236 2790 17389
rect 2916 17236 2982 17389
rect 3108 17236 3174 17389
rect 3300 17236 3356 17389
rect 3784 17236 3850 17389
rect 3976 17236 4042 17389
rect 4168 17236 4234 17389
rect 4360 17236 4426 17389
rect 4552 17236 4618 17389
rect 4744 17236 4810 17389
rect 4936 17236 5002 17389
rect 5128 17236 5184 17389
rect 5612 17236 5678 17389
rect 5804 17236 5870 17389
rect 5996 17236 6062 17389
rect 6188 17236 6254 17389
rect 6380 17236 6446 17389
rect 6572 17236 6638 17389
rect 6764 17236 6830 17389
rect 6956 17236 7012 17389
rect 7440 17236 7506 17389
rect 7632 17236 7698 17389
rect 7824 17236 7890 17389
rect 8016 17236 8082 17389
rect 8208 17236 8274 17389
rect 8400 17236 8466 17389
rect 8592 17236 8658 17389
rect 8784 17236 8840 17389
rect 9268 17236 9334 17389
rect 9460 17236 9526 17389
rect 9652 17236 9718 17389
rect 9844 17236 9910 17389
rect 10036 17236 10102 17389
rect 10228 17236 10294 17389
rect 10420 17236 10486 17389
rect 10612 17236 10668 17389
rect 11096 17236 11162 17389
rect 11288 17236 11354 17389
rect 11480 17236 11546 17389
rect 11672 17236 11738 17389
rect 11864 17236 11930 17389
rect 12056 17236 12122 17389
rect 12248 17236 12314 17389
rect 12440 17236 12496 17389
rect 12924 17236 12990 17389
rect 13116 17236 13182 17389
rect 13308 17236 13374 17389
rect 13500 17236 13566 17389
rect 13692 17236 13758 17389
rect 13884 17236 13950 17389
rect 14076 17236 14142 17389
rect 14268 17236 14324 17389
rect 14752 17236 14818 17389
rect 14944 17236 15010 17389
rect 15136 17236 15202 17389
rect 15328 17236 15394 17389
rect 15520 17236 15586 17389
rect 15712 17236 15778 17389
rect 15904 17236 15970 17389
rect 16096 17236 16152 17389
rect 16580 17236 16646 17389
rect 16772 17236 16838 17389
rect 16964 17236 17030 17389
rect 17156 17236 17222 17389
rect 17348 17236 17414 17389
rect 17540 17236 17606 17389
rect 17732 17236 17798 17389
rect 17924 17236 17980 17389
rect 18408 17236 18474 17389
rect 18600 17236 18666 17389
rect 18792 17236 18858 17389
rect 18984 17236 19050 17389
rect 19176 17236 19242 17389
rect 19368 17236 19434 17389
rect 19560 17236 19626 17389
rect 19752 17236 19808 17389
rect 20236 17236 20302 17389
rect 20428 17236 20494 17389
rect 20620 17236 20686 17389
rect 20812 17236 20878 17389
rect 21004 17236 21070 17389
rect 21196 17236 21262 17389
rect 21388 17236 21454 17389
rect 21580 17236 21636 17389
rect 32 16735 98 16888
rect 224 16735 290 16888
rect 416 16735 482 16888
rect 608 16735 674 16888
rect 800 16735 866 16888
rect 992 16735 1058 16888
rect 1184 16735 1250 16888
rect 1376 16735 1442 16888
rect 1860 16735 1926 16888
rect 2052 16735 2118 16888
rect 2244 16735 2310 16888
rect 2436 16735 2502 16888
rect 2628 16735 2694 16888
rect 2820 16735 2886 16888
rect 3012 16735 3078 16888
rect 3204 16735 3270 16888
rect 3688 16735 3754 16888
rect 3880 16735 3946 16888
rect 4072 16735 4138 16888
rect 4264 16735 4330 16888
rect 4456 16735 4522 16888
rect 4648 16735 4714 16888
rect 4840 16735 4906 16888
rect 5032 16735 5098 16888
rect 5516 16735 5582 16888
rect 5708 16735 5774 16888
rect 5900 16735 5966 16888
rect 6092 16735 6158 16888
rect 6284 16735 6350 16888
rect 6476 16735 6542 16888
rect 6668 16735 6734 16888
rect 6860 16735 6926 16888
rect 7344 16735 7410 16888
rect 7536 16735 7602 16888
rect 7728 16735 7794 16888
rect 7920 16735 7986 16888
rect 8112 16735 8178 16888
rect 8304 16735 8370 16888
rect 8496 16735 8562 16888
rect 8688 16735 8754 16888
rect 9172 16735 9238 16888
rect 9364 16735 9430 16888
rect 9556 16735 9622 16888
rect 9748 16735 9814 16888
rect 9940 16735 10006 16888
rect 10132 16735 10198 16888
rect 10324 16735 10390 16888
rect 10516 16735 10582 16888
rect 11000 16735 11066 16888
rect 11192 16735 11258 16888
rect 11384 16735 11450 16888
rect 11576 16735 11642 16888
rect 11768 16735 11834 16888
rect 11960 16735 12026 16888
rect 12152 16735 12218 16888
rect 12344 16735 12410 16888
rect 12828 16735 12894 16888
rect 13020 16735 13086 16888
rect 13212 16735 13278 16888
rect 13404 16735 13470 16888
rect 13596 16735 13662 16888
rect 13788 16735 13854 16888
rect 13980 16735 14046 16888
rect 14172 16735 14238 16888
rect 14656 16735 14722 16888
rect 14848 16735 14914 16888
rect 15040 16735 15106 16888
rect 15232 16735 15298 16888
rect 15424 16735 15490 16888
rect 15616 16735 15682 16888
rect 15808 16735 15874 16888
rect 16000 16735 16066 16888
rect 16484 16735 16550 16888
rect 16676 16735 16742 16888
rect 16868 16735 16934 16888
rect 17060 16735 17126 16888
rect 17252 16735 17318 16888
rect 17444 16735 17510 16888
rect 17636 16735 17702 16888
rect 17828 16735 17894 16888
rect 18312 16735 18378 16888
rect 18504 16735 18570 16888
rect 18696 16735 18762 16888
rect 18888 16735 18954 16888
rect 19080 16735 19146 16888
rect 19272 16735 19338 16888
rect 19464 16735 19530 16888
rect 19656 16735 19722 16888
rect 20140 16735 20206 16888
rect 20332 16735 20398 16888
rect 20524 16735 20590 16888
rect 20716 16735 20782 16888
rect 20908 16735 20974 16888
rect 21100 16735 21166 16888
rect 21292 16735 21358 16888
rect 21484 16735 21550 16888
rect 128 16522 194 16675
rect 320 16522 386 16675
rect 512 16522 578 16675
rect 704 16522 770 16675
rect 896 16522 962 16675
rect 1088 16522 1154 16675
rect 1280 16522 1346 16675
rect 1472 16522 1528 16675
rect 1956 16522 2022 16675
rect 2148 16522 2214 16675
rect 2340 16522 2406 16675
rect 2532 16522 2598 16675
rect 2724 16522 2790 16675
rect 2916 16522 2982 16675
rect 3108 16522 3174 16675
rect 3300 16522 3356 16675
rect 3784 16522 3850 16675
rect 3976 16522 4042 16675
rect 4168 16522 4234 16675
rect 4360 16522 4426 16675
rect 4552 16522 4618 16675
rect 4744 16522 4810 16675
rect 4936 16522 5002 16675
rect 5128 16522 5184 16675
rect 5612 16522 5678 16675
rect 5804 16522 5870 16675
rect 5996 16522 6062 16675
rect 6188 16522 6254 16675
rect 6380 16522 6446 16675
rect 6572 16522 6638 16675
rect 6764 16522 6830 16675
rect 6956 16522 7012 16675
rect 7440 16522 7506 16675
rect 7632 16522 7698 16675
rect 7824 16522 7890 16675
rect 8016 16522 8082 16675
rect 8208 16522 8274 16675
rect 8400 16522 8466 16675
rect 8592 16522 8658 16675
rect 8784 16522 8840 16675
rect 9268 16522 9334 16675
rect 9460 16522 9526 16675
rect 9652 16522 9718 16675
rect 9844 16522 9910 16675
rect 10036 16522 10102 16675
rect 10228 16522 10294 16675
rect 10420 16522 10486 16675
rect 10612 16522 10668 16675
rect 11096 16522 11162 16675
rect 11288 16522 11354 16675
rect 11480 16522 11546 16675
rect 11672 16522 11738 16675
rect 11864 16522 11930 16675
rect 12056 16522 12122 16675
rect 12248 16522 12314 16675
rect 12440 16522 12496 16675
rect 12924 16522 12990 16675
rect 13116 16522 13182 16675
rect 13308 16522 13374 16675
rect 13500 16522 13566 16675
rect 13692 16522 13758 16675
rect 13884 16522 13950 16675
rect 14076 16522 14142 16675
rect 14268 16522 14324 16675
rect 14752 16522 14818 16675
rect 14944 16522 15010 16675
rect 15136 16522 15202 16675
rect 15328 16522 15394 16675
rect 15520 16522 15586 16675
rect 15712 16522 15778 16675
rect 15904 16522 15970 16675
rect 16096 16522 16152 16675
rect 16580 16522 16646 16675
rect 16772 16522 16838 16675
rect 16964 16522 17030 16675
rect 17156 16522 17222 16675
rect 17348 16522 17414 16675
rect 17540 16522 17606 16675
rect 17732 16522 17798 16675
rect 17924 16522 17980 16675
rect 18408 16522 18474 16675
rect 18600 16522 18666 16675
rect 18792 16522 18858 16675
rect 18984 16522 19050 16675
rect 19176 16522 19242 16675
rect 19368 16522 19434 16675
rect 19560 16522 19626 16675
rect 19752 16522 19808 16675
rect 20236 16522 20302 16675
rect 20428 16522 20494 16675
rect 20620 16522 20686 16675
rect 20812 16522 20878 16675
rect 21004 16522 21070 16675
rect 21196 16522 21262 16675
rect 21388 16522 21454 16675
rect 21580 16522 21636 16675
rect 32 16021 98 16174
rect 224 16021 290 16174
rect 416 16021 482 16174
rect 608 16021 674 16174
rect 800 16021 866 16174
rect 992 16021 1058 16174
rect 1184 16021 1250 16174
rect 1376 16021 1442 16174
rect 1860 16021 1926 16174
rect 2052 16021 2118 16174
rect 2244 16021 2310 16174
rect 2436 16021 2502 16174
rect 2628 16021 2694 16174
rect 2820 16021 2886 16174
rect 3012 16021 3078 16174
rect 3204 16021 3270 16174
rect 3688 16021 3754 16174
rect 3880 16021 3946 16174
rect 4072 16021 4138 16174
rect 4264 16021 4330 16174
rect 4456 16021 4522 16174
rect 4648 16021 4714 16174
rect 4840 16021 4906 16174
rect 5032 16021 5098 16174
rect 5516 16021 5582 16174
rect 5708 16021 5774 16174
rect 5900 16021 5966 16174
rect 6092 16021 6158 16174
rect 6284 16021 6350 16174
rect 6476 16021 6542 16174
rect 6668 16021 6734 16174
rect 6860 16021 6926 16174
rect 7344 16021 7410 16174
rect 7536 16021 7602 16174
rect 7728 16021 7794 16174
rect 7920 16021 7986 16174
rect 8112 16021 8178 16174
rect 8304 16021 8370 16174
rect 8496 16021 8562 16174
rect 8688 16021 8754 16174
rect 9172 16021 9238 16174
rect 9364 16021 9430 16174
rect 9556 16021 9622 16174
rect 9748 16021 9814 16174
rect 9940 16021 10006 16174
rect 10132 16021 10198 16174
rect 10324 16021 10390 16174
rect 10516 16021 10582 16174
rect 11000 16021 11066 16174
rect 11192 16021 11258 16174
rect 11384 16021 11450 16174
rect 11576 16021 11642 16174
rect 11768 16021 11834 16174
rect 11960 16021 12026 16174
rect 12152 16021 12218 16174
rect 12344 16021 12410 16174
rect 12828 16021 12894 16174
rect 13020 16021 13086 16174
rect 13212 16021 13278 16174
rect 13404 16021 13470 16174
rect 13596 16021 13662 16174
rect 13788 16021 13854 16174
rect 13980 16021 14046 16174
rect 14172 16021 14238 16174
rect 14656 16021 14722 16174
rect 14848 16021 14914 16174
rect 15040 16021 15106 16174
rect 15232 16021 15298 16174
rect 15424 16021 15490 16174
rect 15616 16021 15682 16174
rect 15808 16021 15874 16174
rect 16000 16021 16066 16174
rect 16484 16021 16550 16174
rect 16676 16021 16742 16174
rect 16868 16021 16934 16174
rect 17060 16021 17126 16174
rect 17252 16021 17318 16174
rect 17444 16021 17510 16174
rect 17636 16021 17702 16174
rect 17828 16021 17894 16174
rect 18312 16021 18378 16174
rect 18504 16021 18570 16174
rect 18696 16021 18762 16174
rect 18888 16021 18954 16174
rect 19080 16021 19146 16174
rect 19272 16021 19338 16174
rect 19464 16021 19530 16174
rect 19656 16021 19722 16174
rect 20140 16021 20206 16174
rect 20332 16021 20398 16174
rect 20524 16021 20590 16174
rect 20716 16021 20782 16174
rect 20908 16021 20974 16174
rect 21100 16021 21166 16174
rect 21292 16021 21358 16174
rect 21484 16021 21550 16174
rect 128 15808 194 15961
rect 320 15808 386 15961
rect 512 15808 578 15961
rect 704 15808 770 15961
rect 896 15808 962 15961
rect 1088 15808 1154 15961
rect 1280 15808 1346 15961
rect 1472 15808 1528 15961
rect 1956 15808 2022 15961
rect 2148 15808 2214 15961
rect 2340 15808 2406 15961
rect 2532 15808 2598 15961
rect 2724 15808 2790 15961
rect 2916 15808 2982 15961
rect 3108 15808 3174 15961
rect 3300 15808 3356 15961
rect 3784 15808 3850 15961
rect 3976 15808 4042 15961
rect 4168 15808 4234 15961
rect 4360 15808 4426 15961
rect 4552 15808 4618 15961
rect 4744 15808 4810 15961
rect 4936 15808 5002 15961
rect 5128 15808 5184 15961
rect 5612 15808 5678 15961
rect 5804 15808 5870 15961
rect 5996 15808 6062 15961
rect 6188 15808 6254 15961
rect 6380 15808 6446 15961
rect 6572 15808 6638 15961
rect 6764 15808 6830 15961
rect 6956 15808 7012 15961
rect 7440 15808 7506 15961
rect 7632 15808 7698 15961
rect 7824 15808 7890 15961
rect 8016 15808 8082 15961
rect 8208 15808 8274 15961
rect 8400 15808 8466 15961
rect 8592 15808 8658 15961
rect 8784 15808 8840 15961
rect 9268 15808 9334 15961
rect 9460 15808 9526 15961
rect 9652 15808 9718 15961
rect 9844 15808 9910 15961
rect 10036 15808 10102 15961
rect 10228 15808 10294 15961
rect 10420 15808 10486 15961
rect 10612 15808 10668 15961
rect 11096 15808 11162 15961
rect 11288 15808 11354 15961
rect 11480 15808 11546 15961
rect 11672 15808 11738 15961
rect 11864 15808 11930 15961
rect 12056 15808 12122 15961
rect 12248 15808 12314 15961
rect 12440 15808 12496 15961
rect 12924 15808 12990 15961
rect 13116 15808 13182 15961
rect 13308 15808 13374 15961
rect 13500 15808 13566 15961
rect 13692 15808 13758 15961
rect 13884 15808 13950 15961
rect 14076 15808 14142 15961
rect 14268 15808 14324 15961
rect 14752 15808 14818 15961
rect 14944 15808 15010 15961
rect 15136 15808 15202 15961
rect 15328 15808 15394 15961
rect 15520 15808 15586 15961
rect 15712 15808 15778 15961
rect 15904 15808 15970 15961
rect 16096 15808 16152 15961
rect 16580 15808 16646 15961
rect 16772 15808 16838 15961
rect 16964 15808 17030 15961
rect 17156 15808 17222 15961
rect 17348 15808 17414 15961
rect 17540 15808 17606 15961
rect 17732 15808 17798 15961
rect 17924 15808 17980 15961
rect 18408 15808 18474 15961
rect 18600 15808 18666 15961
rect 18792 15808 18858 15961
rect 18984 15808 19050 15961
rect 19176 15808 19242 15961
rect 19368 15808 19434 15961
rect 19560 15808 19626 15961
rect 19752 15808 19808 15961
rect 20236 15808 20302 15961
rect 20428 15808 20494 15961
rect 20620 15808 20686 15961
rect 20812 15808 20878 15961
rect 21004 15808 21070 15961
rect 21196 15808 21262 15961
rect 21388 15808 21454 15961
rect 21580 15808 21636 15961
rect 32 15307 98 15460
rect 224 15307 290 15460
rect 416 15307 482 15460
rect 608 15307 674 15460
rect 800 15307 866 15460
rect 992 15307 1058 15460
rect 1184 15307 1250 15460
rect 1376 15307 1442 15460
rect 1860 15307 1926 15460
rect 2052 15307 2118 15460
rect 2244 15307 2310 15460
rect 2436 15307 2502 15460
rect 2628 15307 2694 15460
rect 2820 15307 2886 15460
rect 3012 15307 3078 15460
rect 3204 15307 3270 15460
rect 3688 15307 3754 15460
rect 3880 15307 3946 15460
rect 4072 15307 4138 15460
rect 4264 15307 4330 15460
rect 4456 15307 4522 15460
rect 4648 15307 4714 15460
rect 4840 15307 4906 15460
rect 5032 15307 5098 15460
rect 5516 15307 5582 15460
rect 5708 15307 5774 15460
rect 5900 15307 5966 15460
rect 6092 15307 6158 15460
rect 6284 15307 6350 15460
rect 6476 15307 6542 15460
rect 6668 15307 6734 15460
rect 6860 15307 6926 15460
rect 7344 15307 7410 15460
rect 7536 15307 7602 15460
rect 7728 15307 7794 15460
rect 7920 15307 7986 15460
rect 8112 15307 8178 15460
rect 8304 15307 8370 15460
rect 8496 15307 8562 15460
rect 8688 15307 8754 15460
rect 9172 15307 9238 15460
rect 9364 15307 9430 15460
rect 9556 15307 9622 15460
rect 9748 15307 9814 15460
rect 9940 15307 10006 15460
rect 10132 15307 10198 15460
rect 10324 15307 10390 15460
rect 10516 15307 10582 15460
rect 11000 15307 11066 15460
rect 11192 15307 11258 15460
rect 11384 15307 11450 15460
rect 11576 15307 11642 15460
rect 11768 15307 11834 15460
rect 11960 15307 12026 15460
rect 12152 15307 12218 15460
rect 12344 15307 12410 15460
rect 12828 15307 12894 15460
rect 13020 15307 13086 15460
rect 13212 15307 13278 15460
rect 13404 15307 13470 15460
rect 13596 15307 13662 15460
rect 13788 15307 13854 15460
rect 13980 15307 14046 15460
rect 14172 15307 14238 15460
rect 14656 15307 14722 15460
rect 14848 15307 14914 15460
rect 15040 15307 15106 15460
rect 15232 15307 15298 15460
rect 15424 15307 15490 15460
rect 15616 15307 15682 15460
rect 15808 15307 15874 15460
rect 16000 15307 16066 15460
rect 16484 15307 16550 15460
rect 16676 15307 16742 15460
rect 16868 15307 16934 15460
rect 17060 15307 17126 15460
rect 17252 15307 17318 15460
rect 17444 15307 17510 15460
rect 17636 15307 17702 15460
rect 17828 15307 17894 15460
rect 18312 15307 18378 15460
rect 18504 15307 18570 15460
rect 18696 15307 18762 15460
rect 18888 15307 18954 15460
rect 19080 15307 19146 15460
rect 19272 15307 19338 15460
rect 19464 15307 19530 15460
rect 19656 15307 19722 15460
rect 20140 15307 20206 15460
rect 20332 15307 20398 15460
rect 20524 15307 20590 15460
rect 20716 15307 20782 15460
rect 20908 15307 20974 15460
rect 21100 15307 21166 15460
rect 21292 15307 21358 15460
rect 21484 15307 21550 15460
rect 128 15094 194 15247
rect 320 15094 386 15247
rect 512 15094 578 15247
rect 704 15094 770 15247
rect 896 15094 962 15247
rect 1088 15094 1154 15247
rect 1280 15094 1346 15247
rect 1472 15094 1528 15247
rect 1956 15094 2022 15247
rect 2148 15094 2214 15247
rect 2340 15094 2406 15247
rect 2532 15094 2598 15247
rect 2724 15094 2790 15247
rect 2916 15094 2982 15247
rect 3108 15094 3174 15247
rect 3300 15094 3356 15247
rect 3784 15094 3850 15247
rect 3976 15094 4042 15247
rect 4168 15094 4234 15247
rect 4360 15094 4426 15247
rect 4552 15094 4618 15247
rect 4744 15094 4810 15247
rect 4936 15094 5002 15247
rect 5128 15094 5184 15247
rect 5612 15094 5678 15247
rect 5804 15094 5870 15247
rect 5996 15094 6062 15247
rect 6188 15094 6254 15247
rect 6380 15094 6446 15247
rect 6572 15094 6638 15247
rect 6764 15094 6830 15247
rect 6956 15094 7012 15247
rect 7440 15094 7506 15247
rect 7632 15094 7698 15247
rect 7824 15094 7890 15247
rect 8016 15094 8082 15247
rect 8208 15094 8274 15247
rect 8400 15094 8466 15247
rect 8592 15094 8658 15247
rect 8784 15094 8840 15247
rect 9268 15094 9334 15247
rect 9460 15094 9526 15247
rect 9652 15094 9718 15247
rect 9844 15094 9910 15247
rect 10036 15094 10102 15247
rect 10228 15094 10294 15247
rect 10420 15094 10486 15247
rect 10612 15094 10668 15247
rect 11096 15094 11162 15247
rect 11288 15094 11354 15247
rect 11480 15094 11546 15247
rect 11672 15094 11738 15247
rect 11864 15094 11930 15247
rect 12056 15094 12122 15247
rect 12248 15094 12314 15247
rect 12440 15094 12496 15247
rect 12924 15094 12990 15247
rect 13116 15094 13182 15247
rect 13308 15094 13374 15247
rect 13500 15094 13566 15247
rect 13692 15094 13758 15247
rect 13884 15094 13950 15247
rect 14076 15094 14142 15247
rect 14268 15094 14324 15247
rect 14752 15094 14818 15247
rect 14944 15094 15010 15247
rect 15136 15094 15202 15247
rect 15328 15094 15394 15247
rect 15520 15094 15586 15247
rect 15712 15094 15778 15247
rect 15904 15094 15970 15247
rect 16096 15094 16152 15247
rect 16580 15094 16646 15247
rect 16772 15094 16838 15247
rect 16964 15094 17030 15247
rect 17156 15094 17222 15247
rect 17348 15094 17414 15247
rect 17540 15094 17606 15247
rect 17732 15094 17798 15247
rect 17924 15094 17980 15247
rect 18408 15094 18474 15247
rect 18600 15094 18666 15247
rect 18792 15094 18858 15247
rect 18984 15094 19050 15247
rect 19176 15094 19242 15247
rect 19368 15094 19434 15247
rect 19560 15094 19626 15247
rect 19752 15094 19808 15247
rect 20236 15094 20302 15247
rect 20428 15094 20494 15247
rect 20620 15094 20686 15247
rect 20812 15094 20878 15247
rect 21004 15094 21070 15247
rect 21196 15094 21262 15247
rect 21388 15094 21454 15247
rect 21580 15094 21636 15247
rect 32 14593 98 14746
rect 224 14593 290 14746
rect 416 14593 482 14746
rect 608 14593 674 14746
rect 800 14593 866 14746
rect 992 14593 1058 14746
rect 1184 14593 1250 14746
rect 1376 14593 1442 14746
rect 1860 14593 1926 14746
rect 2052 14593 2118 14746
rect 2244 14593 2310 14746
rect 2436 14593 2502 14746
rect 2628 14593 2694 14746
rect 2820 14593 2886 14746
rect 3012 14593 3078 14746
rect 3204 14593 3270 14746
rect 3688 14593 3754 14746
rect 3880 14593 3946 14746
rect 4072 14593 4138 14746
rect 4264 14593 4330 14746
rect 4456 14593 4522 14746
rect 4648 14593 4714 14746
rect 4840 14593 4906 14746
rect 5032 14593 5098 14746
rect 5516 14593 5582 14746
rect 5708 14593 5774 14746
rect 5900 14593 5966 14746
rect 6092 14593 6158 14746
rect 6284 14593 6350 14746
rect 6476 14593 6542 14746
rect 6668 14593 6734 14746
rect 6860 14593 6926 14746
rect 7344 14593 7410 14746
rect 7536 14593 7602 14746
rect 7728 14593 7794 14746
rect 7920 14593 7986 14746
rect 8112 14593 8178 14746
rect 8304 14593 8370 14746
rect 8496 14593 8562 14746
rect 8688 14593 8754 14746
rect 9172 14593 9238 14746
rect 9364 14593 9430 14746
rect 9556 14593 9622 14746
rect 9748 14593 9814 14746
rect 9940 14593 10006 14746
rect 10132 14593 10198 14746
rect 10324 14593 10390 14746
rect 10516 14593 10582 14746
rect 11000 14593 11066 14746
rect 11192 14593 11258 14746
rect 11384 14593 11450 14746
rect 11576 14593 11642 14746
rect 11768 14593 11834 14746
rect 11960 14593 12026 14746
rect 12152 14593 12218 14746
rect 12344 14593 12410 14746
rect 12828 14593 12894 14746
rect 13020 14593 13086 14746
rect 13212 14593 13278 14746
rect 13404 14593 13470 14746
rect 13596 14593 13662 14746
rect 13788 14593 13854 14746
rect 13980 14593 14046 14746
rect 14172 14593 14238 14746
rect 14656 14593 14722 14746
rect 14848 14593 14914 14746
rect 15040 14593 15106 14746
rect 15232 14593 15298 14746
rect 15424 14593 15490 14746
rect 15616 14593 15682 14746
rect 15808 14593 15874 14746
rect 16000 14593 16066 14746
rect 16484 14593 16550 14746
rect 16676 14593 16742 14746
rect 16868 14593 16934 14746
rect 17060 14593 17126 14746
rect 17252 14593 17318 14746
rect 17444 14593 17510 14746
rect 17636 14593 17702 14746
rect 17828 14593 17894 14746
rect 18312 14593 18378 14746
rect 18504 14593 18570 14746
rect 18696 14593 18762 14746
rect 18888 14593 18954 14746
rect 19080 14593 19146 14746
rect 19272 14593 19338 14746
rect 19464 14593 19530 14746
rect 19656 14593 19722 14746
rect 20140 14593 20206 14746
rect 20332 14593 20398 14746
rect 20524 14593 20590 14746
rect 20716 14593 20782 14746
rect 20908 14593 20974 14746
rect 21100 14593 21166 14746
rect 21292 14593 21358 14746
rect 21484 14593 21550 14746
rect 128 14380 194 14533
rect 320 14380 386 14533
rect 512 14380 578 14533
rect 704 14380 770 14533
rect 896 14380 962 14533
rect 1088 14380 1154 14533
rect 1280 14380 1346 14533
rect 1472 14380 1528 14533
rect 1956 14380 2022 14533
rect 2148 14380 2214 14533
rect 2340 14380 2406 14533
rect 2532 14380 2598 14533
rect 2724 14380 2790 14533
rect 2916 14380 2982 14533
rect 3108 14380 3174 14533
rect 3300 14380 3356 14533
rect 3784 14380 3850 14533
rect 3976 14380 4042 14533
rect 4168 14380 4234 14533
rect 4360 14380 4426 14533
rect 4552 14380 4618 14533
rect 4744 14380 4810 14533
rect 4936 14380 5002 14533
rect 5128 14380 5184 14533
rect 5612 14380 5678 14533
rect 5804 14380 5870 14533
rect 5996 14380 6062 14533
rect 6188 14380 6254 14533
rect 6380 14380 6446 14533
rect 6572 14380 6638 14533
rect 6764 14380 6830 14533
rect 6956 14380 7012 14533
rect 7440 14380 7506 14533
rect 7632 14380 7698 14533
rect 7824 14380 7890 14533
rect 8016 14380 8082 14533
rect 8208 14380 8274 14533
rect 8400 14380 8466 14533
rect 8592 14380 8658 14533
rect 8784 14380 8840 14533
rect 9268 14380 9334 14533
rect 9460 14380 9526 14533
rect 9652 14380 9718 14533
rect 9844 14380 9910 14533
rect 10036 14380 10102 14533
rect 10228 14380 10294 14533
rect 10420 14380 10486 14533
rect 10612 14380 10668 14533
rect 11096 14380 11162 14533
rect 11288 14380 11354 14533
rect 11480 14380 11546 14533
rect 11672 14380 11738 14533
rect 11864 14380 11930 14533
rect 12056 14380 12122 14533
rect 12248 14380 12314 14533
rect 12440 14380 12496 14533
rect 12924 14380 12990 14533
rect 13116 14380 13182 14533
rect 13308 14380 13374 14533
rect 13500 14380 13566 14533
rect 13692 14380 13758 14533
rect 13884 14380 13950 14533
rect 14076 14380 14142 14533
rect 14268 14380 14324 14533
rect 14752 14380 14818 14533
rect 14944 14380 15010 14533
rect 15136 14380 15202 14533
rect 15328 14380 15394 14533
rect 15520 14380 15586 14533
rect 15712 14380 15778 14533
rect 15904 14380 15970 14533
rect 16096 14380 16152 14533
rect 16580 14380 16646 14533
rect 16772 14380 16838 14533
rect 16964 14380 17030 14533
rect 17156 14380 17222 14533
rect 17348 14380 17414 14533
rect 17540 14380 17606 14533
rect 17732 14380 17798 14533
rect 17924 14380 17980 14533
rect 18408 14380 18474 14533
rect 18600 14380 18666 14533
rect 18792 14380 18858 14533
rect 18984 14380 19050 14533
rect 19176 14380 19242 14533
rect 19368 14380 19434 14533
rect 19560 14380 19626 14533
rect 19752 14380 19808 14533
rect 20236 14380 20302 14533
rect 20428 14380 20494 14533
rect 20620 14380 20686 14533
rect 20812 14380 20878 14533
rect 21004 14380 21070 14533
rect 21196 14380 21262 14533
rect 21388 14380 21454 14533
rect 21580 14380 21636 14533
rect 32 13879 98 14032
rect 224 13879 290 14032
rect 416 13879 482 14032
rect 608 13879 674 14032
rect 800 13879 866 14032
rect 992 13879 1058 14032
rect 1184 13879 1250 14032
rect 1376 13879 1442 14032
rect 1860 13879 1926 14032
rect 2052 13879 2118 14032
rect 2244 13879 2310 14032
rect 2436 13879 2502 14032
rect 2628 13879 2694 14032
rect 2820 13879 2886 14032
rect 3012 13879 3078 14032
rect 3204 13879 3270 14032
rect 3688 13879 3754 14032
rect 3880 13879 3946 14032
rect 4072 13879 4138 14032
rect 4264 13879 4330 14032
rect 4456 13879 4522 14032
rect 4648 13879 4714 14032
rect 4840 13879 4906 14032
rect 5032 13879 5098 14032
rect 5516 13879 5582 14032
rect 5708 13879 5774 14032
rect 5900 13879 5966 14032
rect 6092 13879 6158 14032
rect 6284 13879 6350 14032
rect 6476 13879 6542 14032
rect 6668 13879 6734 14032
rect 6860 13879 6926 14032
rect 7344 13879 7410 14032
rect 7536 13879 7602 14032
rect 7728 13879 7794 14032
rect 7920 13879 7986 14032
rect 8112 13879 8178 14032
rect 8304 13879 8370 14032
rect 8496 13879 8562 14032
rect 8688 13879 8754 14032
rect 9172 13879 9238 14032
rect 9364 13879 9430 14032
rect 9556 13879 9622 14032
rect 9748 13879 9814 14032
rect 9940 13879 10006 14032
rect 10132 13879 10198 14032
rect 10324 13879 10390 14032
rect 10516 13879 10582 14032
rect 11000 13879 11066 14032
rect 11192 13879 11258 14032
rect 11384 13879 11450 14032
rect 11576 13879 11642 14032
rect 11768 13879 11834 14032
rect 11960 13879 12026 14032
rect 12152 13879 12218 14032
rect 12344 13879 12410 14032
rect 12828 13879 12894 14032
rect 13020 13879 13086 14032
rect 13212 13879 13278 14032
rect 13404 13879 13470 14032
rect 13596 13879 13662 14032
rect 13788 13879 13854 14032
rect 13980 13879 14046 14032
rect 14172 13879 14238 14032
rect 14656 13879 14722 14032
rect 14848 13879 14914 14032
rect 15040 13879 15106 14032
rect 15232 13879 15298 14032
rect 15424 13879 15490 14032
rect 15616 13879 15682 14032
rect 15808 13879 15874 14032
rect 16000 13879 16066 14032
rect 16484 13879 16550 14032
rect 16676 13879 16742 14032
rect 16868 13879 16934 14032
rect 17060 13879 17126 14032
rect 17252 13879 17318 14032
rect 17444 13879 17510 14032
rect 17636 13879 17702 14032
rect 17828 13879 17894 14032
rect 18312 13879 18378 14032
rect 18504 13879 18570 14032
rect 18696 13879 18762 14032
rect 18888 13879 18954 14032
rect 19080 13879 19146 14032
rect 19272 13879 19338 14032
rect 19464 13879 19530 14032
rect 19656 13879 19722 14032
rect 20140 13879 20206 14032
rect 20332 13879 20398 14032
rect 20524 13879 20590 14032
rect 20716 13879 20782 14032
rect 20908 13879 20974 14032
rect 21100 13879 21166 14032
rect 21292 13879 21358 14032
rect 21484 13879 21550 14032
rect 128 13666 194 13819
rect 320 13666 386 13819
rect 512 13666 578 13819
rect 704 13666 770 13819
rect 896 13666 962 13819
rect 1088 13666 1154 13819
rect 1280 13666 1346 13819
rect 1472 13666 1528 13819
rect 1956 13666 2022 13819
rect 2148 13666 2214 13819
rect 2340 13666 2406 13819
rect 2532 13666 2598 13819
rect 2724 13666 2790 13819
rect 2916 13666 2982 13819
rect 3108 13666 3174 13819
rect 3300 13666 3356 13819
rect 3784 13666 3850 13819
rect 3976 13666 4042 13819
rect 4168 13666 4234 13819
rect 4360 13666 4426 13819
rect 4552 13666 4618 13819
rect 4744 13666 4810 13819
rect 4936 13666 5002 13819
rect 5128 13666 5184 13819
rect 5612 13666 5678 13819
rect 5804 13666 5870 13819
rect 5996 13666 6062 13819
rect 6188 13666 6254 13819
rect 6380 13666 6446 13819
rect 6572 13666 6638 13819
rect 6764 13666 6830 13819
rect 6956 13666 7012 13819
rect 7440 13666 7506 13819
rect 7632 13666 7698 13819
rect 7824 13666 7890 13819
rect 8016 13666 8082 13819
rect 8208 13666 8274 13819
rect 8400 13666 8466 13819
rect 8592 13666 8658 13819
rect 8784 13666 8840 13819
rect 9268 13666 9334 13819
rect 9460 13666 9526 13819
rect 9652 13666 9718 13819
rect 9844 13666 9910 13819
rect 10036 13666 10102 13819
rect 10228 13666 10294 13819
rect 10420 13666 10486 13819
rect 10612 13666 10668 13819
rect 11096 13666 11162 13819
rect 11288 13666 11354 13819
rect 11480 13666 11546 13819
rect 11672 13666 11738 13819
rect 11864 13666 11930 13819
rect 12056 13666 12122 13819
rect 12248 13666 12314 13819
rect 12440 13666 12496 13819
rect 12924 13666 12990 13819
rect 13116 13666 13182 13819
rect 13308 13666 13374 13819
rect 13500 13666 13566 13819
rect 13692 13666 13758 13819
rect 13884 13666 13950 13819
rect 14076 13666 14142 13819
rect 14268 13666 14324 13819
rect 14752 13666 14818 13819
rect 14944 13666 15010 13819
rect 15136 13666 15202 13819
rect 15328 13666 15394 13819
rect 15520 13666 15586 13819
rect 15712 13666 15778 13819
rect 15904 13666 15970 13819
rect 16096 13666 16152 13819
rect 16580 13666 16646 13819
rect 16772 13666 16838 13819
rect 16964 13666 17030 13819
rect 17156 13666 17222 13819
rect 17348 13666 17414 13819
rect 17540 13666 17606 13819
rect 17732 13666 17798 13819
rect 17924 13666 17980 13819
rect 18408 13666 18474 13819
rect 18600 13666 18666 13819
rect 18792 13666 18858 13819
rect 18984 13666 19050 13819
rect 19176 13666 19242 13819
rect 19368 13666 19434 13819
rect 19560 13666 19626 13819
rect 19752 13666 19808 13819
rect 20236 13666 20302 13819
rect 20428 13666 20494 13819
rect 20620 13666 20686 13819
rect 20812 13666 20878 13819
rect 21004 13666 21070 13819
rect 21196 13666 21262 13819
rect 21388 13666 21454 13819
rect 21580 13666 21636 13819
rect 32 13165 98 13318
rect 224 13165 290 13318
rect 416 13165 482 13318
rect 608 13165 674 13318
rect 800 13165 866 13318
rect 992 13165 1058 13318
rect 1184 13165 1250 13318
rect 1376 13165 1442 13318
rect 1860 13165 1926 13318
rect 2052 13165 2118 13318
rect 2244 13165 2310 13318
rect 2436 13165 2502 13318
rect 2628 13165 2694 13318
rect 2820 13165 2886 13318
rect 3012 13165 3078 13318
rect 3204 13165 3270 13318
rect 3688 13165 3754 13318
rect 3880 13165 3946 13318
rect 4072 13165 4138 13318
rect 4264 13165 4330 13318
rect 4456 13165 4522 13318
rect 4648 13165 4714 13318
rect 4840 13165 4906 13318
rect 5032 13165 5098 13318
rect 5516 13165 5582 13318
rect 5708 13165 5774 13318
rect 5900 13165 5966 13318
rect 6092 13165 6158 13318
rect 6284 13165 6350 13318
rect 6476 13165 6542 13318
rect 6668 13165 6734 13318
rect 6860 13165 6926 13318
rect 7344 13165 7410 13318
rect 7536 13165 7602 13318
rect 7728 13165 7794 13318
rect 7920 13165 7986 13318
rect 8112 13165 8178 13318
rect 8304 13165 8370 13318
rect 8496 13165 8562 13318
rect 8688 13165 8754 13318
rect 9172 13165 9238 13318
rect 9364 13165 9430 13318
rect 9556 13165 9622 13318
rect 9748 13165 9814 13318
rect 9940 13165 10006 13318
rect 10132 13165 10198 13318
rect 10324 13165 10390 13318
rect 10516 13165 10582 13318
rect 11000 13165 11066 13318
rect 11192 13165 11258 13318
rect 11384 13165 11450 13318
rect 11576 13165 11642 13318
rect 11768 13165 11834 13318
rect 11960 13165 12026 13318
rect 12152 13165 12218 13318
rect 12344 13165 12410 13318
rect 12828 13165 12894 13318
rect 13020 13165 13086 13318
rect 13212 13165 13278 13318
rect 13404 13165 13470 13318
rect 13596 13165 13662 13318
rect 13788 13165 13854 13318
rect 13980 13165 14046 13318
rect 14172 13165 14238 13318
rect 14656 13165 14722 13318
rect 14848 13165 14914 13318
rect 15040 13165 15106 13318
rect 15232 13165 15298 13318
rect 15424 13165 15490 13318
rect 15616 13165 15682 13318
rect 15808 13165 15874 13318
rect 16000 13165 16066 13318
rect 16484 13165 16550 13318
rect 16676 13165 16742 13318
rect 16868 13165 16934 13318
rect 17060 13165 17126 13318
rect 17252 13165 17318 13318
rect 17444 13165 17510 13318
rect 17636 13165 17702 13318
rect 17828 13165 17894 13318
rect 18312 13165 18378 13318
rect 18504 13165 18570 13318
rect 18696 13165 18762 13318
rect 18888 13165 18954 13318
rect 19080 13165 19146 13318
rect 19272 13165 19338 13318
rect 19464 13165 19530 13318
rect 19656 13165 19722 13318
rect 20140 13165 20206 13318
rect 20332 13165 20398 13318
rect 20524 13165 20590 13318
rect 20716 13165 20782 13318
rect 20908 13165 20974 13318
rect 21100 13165 21166 13318
rect 21292 13165 21358 13318
rect 21484 13165 21550 13318
rect 128 12952 194 13105
rect 320 12952 386 13105
rect 512 12952 578 13105
rect 704 12952 770 13105
rect 896 12952 962 13105
rect 1088 12952 1154 13105
rect 1280 12952 1346 13105
rect 1472 12952 1528 13105
rect 1956 12952 2022 13105
rect 2148 12952 2214 13105
rect 2340 12952 2406 13105
rect 2532 12952 2598 13105
rect 2724 12952 2790 13105
rect 2916 12952 2982 13105
rect 3108 12952 3174 13105
rect 3300 12952 3356 13105
rect 3784 12952 3850 13105
rect 3976 12952 4042 13105
rect 4168 12952 4234 13105
rect 4360 12952 4426 13105
rect 4552 12952 4618 13105
rect 4744 12952 4810 13105
rect 4936 12952 5002 13105
rect 5128 12952 5184 13105
rect 5612 12952 5678 13105
rect 5804 12952 5870 13105
rect 5996 12952 6062 13105
rect 6188 12952 6254 13105
rect 6380 12952 6446 13105
rect 6572 12952 6638 13105
rect 6764 12952 6830 13105
rect 6956 12952 7012 13105
rect 7440 12952 7506 13105
rect 7632 12952 7698 13105
rect 7824 12952 7890 13105
rect 8016 12952 8082 13105
rect 8208 12952 8274 13105
rect 8400 12952 8466 13105
rect 8592 12952 8658 13105
rect 8784 12952 8840 13105
rect 9268 12952 9334 13105
rect 9460 12952 9526 13105
rect 9652 12952 9718 13105
rect 9844 12952 9910 13105
rect 10036 12952 10102 13105
rect 10228 12952 10294 13105
rect 10420 12952 10486 13105
rect 10612 12952 10668 13105
rect 11096 12952 11162 13105
rect 11288 12952 11354 13105
rect 11480 12952 11546 13105
rect 11672 12952 11738 13105
rect 11864 12952 11930 13105
rect 12056 12952 12122 13105
rect 12248 12952 12314 13105
rect 12440 12952 12496 13105
rect 12924 12952 12990 13105
rect 13116 12952 13182 13105
rect 13308 12952 13374 13105
rect 13500 12952 13566 13105
rect 13692 12952 13758 13105
rect 13884 12952 13950 13105
rect 14076 12952 14142 13105
rect 14268 12952 14324 13105
rect 14752 12952 14818 13105
rect 14944 12952 15010 13105
rect 15136 12952 15202 13105
rect 15328 12952 15394 13105
rect 15520 12952 15586 13105
rect 15712 12952 15778 13105
rect 15904 12952 15970 13105
rect 16096 12952 16152 13105
rect 16580 12952 16646 13105
rect 16772 12952 16838 13105
rect 16964 12952 17030 13105
rect 17156 12952 17222 13105
rect 17348 12952 17414 13105
rect 17540 12952 17606 13105
rect 17732 12952 17798 13105
rect 17924 12952 17980 13105
rect 18408 12952 18474 13105
rect 18600 12952 18666 13105
rect 18792 12952 18858 13105
rect 18984 12952 19050 13105
rect 19176 12952 19242 13105
rect 19368 12952 19434 13105
rect 19560 12952 19626 13105
rect 19752 12952 19808 13105
rect 20236 12952 20302 13105
rect 20428 12952 20494 13105
rect 20620 12952 20686 13105
rect 20812 12952 20878 13105
rect 21004 12952 21070 13105
rect 21196 12952 21262 13105
rect 21388 12952 21454 13105
rect 21580 12952 21636 13105
rect 32 12451 98 12604
rect 224 12451 290 12604
rect 416 12451 482 12604
rect 608 12451 674 12604
rect 800 12451 866 12604
rect 992 12451 1058 12604
rect 1184 12451 1250 12604
rect 1376 12451 1442 12604
rect 1860 12451 1926 12604
rect 2052 12451 2118 12604
rect 2244 12451 2310 12604
rect 2436 12451 2502 12604
rect 2628 12451 2694 12604
rect 2820 12451 2886 12604
rect 3012 12451 3078 12604
rect 3204 12451 3270 12604
rect 3688 12451 3754 12604
rect 3880 12451 3946 12604
rect 4072 12451 4138 12604
rect 4264 12451 4330 12604
rect 4456 12451 4522 12604
rect 4648 12451 4714 12604
rect 4840 12451 4906 12604
rect 5032 12451 5098 12604
rect 5516 12451 5582 12604
rect 5708 12451 5774 12604
rect 5900 12451 5966 12604
rect 6092 12451 6158 12604
rect 6284 12451 6350 12604
rect 6476 12451 6542 12604
rect 6668 12451 6734 12604
rect 6860 12451 6926 12604
rect 7344 12451 7410 12604
rect 7536 12451 7602 12604
rect 7728 12451 7794 12604
rect 7920 12451 7986 12604
rect 8112 12451 8178 12604
rect 8304 12451 8370 12604
rect 8496 12451 8562 12604
rect 8688 12451 8754 12604
rect 9172 12451 9238 12604
rect 9364 12451 9430 12604
rect 9556 12451 9622 12604
rect 9748 12451 9814 12604
rect 9940 12451 10006 12604
rect 10132 12451 10198 12604
rect 10324 12451 10390 12604
rect 10516 12451 10582 12604
rect 11000 12451 11066 12604
rect 11192 12451 11258 12604
rect 11384 12451 11450 12604
rect 11576 12451 11642 12604
rect 11768 12451 11834 12604
rect 11960 12451 12026 12604
rect 12152 12451 12218 12604
rect 12344 12451 12410 12604
rect 12828 12451 12894 12604
rect 13020 12451 13086 12604
rect 13212 12451 13278 12604
rect 13404 12451 13470 12604
rect 13596 12451 13662 12604
rect 13788 12451 13854 12604
rect 13980 12451 14046 12604
rect 14172 12451 14238 12604
rect 14656 12451 14722 12604
rect 14848 12451 14914 12604
rect 15040 12451 15106 12604
rect 15232 12451 15298 12604
rect 15424 12451 15490 12604
rect 15616 12451 15682 12604
rect 15808 12451 15874 12604
rect 16000 12451 16066 12604
rect 16484 12451 16550 12604
rect 16676 12451 16742 12604
rect 16868 12451 16934 12604
rect 17060 12451 17126 12604
rect 17252 12451 17318 12604
rect 17444 12451 17510 12604
rect 17636 12451 17702 12604
rect 17828 12451 17894 12604
rect 18312 12451 18378 12604
rect 18504 12451 18570 12604
rect 18696 12451 18762 12604
rect 18888 12451 18954 12604
rect 19080 12451 19146 12604
rect 19272 12451 19338 12604
rect 19464 12451 19530 12604
rect 19656 12451 19722 12604
rect 20140 12451 20206 12604
rect 20332 12451 20398 12604
rect 20524 12451 20590 12604
rect 20716 12451 20782 12604
rect 20908 12451 20974 12604
rect 21100 12451 21166 12604
rect 21292 12451 21358 12604
rect 21484 12451 21550 12604
rect 128 12238 194 12391
rect 320 12238 386 12391
rect 512 12238 578 12391
rect 704 12238 770 12391
rect 896 12238 962 12391
rect 1088 12238 1154 12391
rect 1280 12238 1346 12391
rect 1472 12238 1528 12391
rect 1956 12238 2022 12391
rect 2148 12238 2214 12391
rect 2340 12238 2406 12391
rect 2532 12238 2598 12391
rect 2724 12238 2790 12391
rect 2916 12238 2982 12391
rect 3108 12238 3174 12391
rect 3300 12238 3356 12391
rect 3784 12238 3850 12391
rect 3976 12238 4042 12391
rect 4168 12238 4234 12391
rect 4360 12238 4426 12391
rect 4552 12238 4618 12391
rect 4744 12238 4810 12391
rect 4936 12238 5002 12391
rect 5128 12238 5184 12391
rect 5612 12238 5678 12391
rect 5804 12238 5870 12391
rect 5996 12238 6062 12391
rect 6188 12238 6254 12391
rect 6380 12238 6446 12391
rect 6572 12238 6638 12391
rect 6764 12238 6830 12391
rect 6956 12238 7012 12391
rect 7440 12238 7506 12391
rect 7632 12238 7698 12391
rect 7824 12238 7890 12391
rect 8016 12238 8082 12391
rect 8208 12238 8274 12391
rect 8400 12238 8466 12391
rect 8592 12238 8658 12391
rect 8784 12238 8840 12391
rect 9268 12238 9334 12391
rect 9460 12238 9526 12391
rect 9652 12238 9718 12391
rect 9844 12238 9910 12391
rect 10036 12238 10102 12391
rect 10228 12238 10294 12391
rect 10420 12238 10486 12391
rect 10612 12238 10668 12391
rect 11096 12238 11162 12391
rect 11288 12238 11354 12391
rect 11480 12238 11546 12391
rect 11672 12238 11738 12391
rect 11864 12238 11930 12391
rect 12056 12238 12122 12391
rect 12248 12238 12314 12391
rect 12440 12238 12496 12391
rect 12924 12238 12990 12391
rect 13116 12238 13182 12391
rect 13308 12238 13374 12391
rect 13500 12238 13566 12391
rect 13692 12238 13758 12391
rect 13884 12238 13950 12391
rect 14076 12238 14142 12391
rect 14268 12238 14324 12391
rect 14752 12238 14818 12391
rect 14944 12238 15010 12391
rect 15136 12238 15202 12391
rect 15328 12238 15394 12391
rect 15520 12238 15586 12391
rect 15712 12238 15778 12391
rect 15904 12238 15970 12391
rect 16096 12238 16152 12391
rect 16580 12238 16646 12391
rect 16772 12238 16838 12391
rect 16964 12238 17030 12391
rect 17156 12238 17222 12391
rect 17348 12238 17414 12391
rect 17540 12238 17606 12391
rect 17732 12238 17798 12391
rect 17924 12238 17980 12391
rect 18408 12238 18474 12391
rect 18600 12238 18666 12391
rect 18792 12238 18858 12391
rect 18984 12238 19050 12391
rect 19176 12238 19242 12391
rect 19368 12238 19434 12391
rect 19560 12238 19626 12391
rect 19752 12238 19808 12391
rect 20236 12238 20302 12391
rect 20428 12238 20494 12391
rect 20620 12238 20686 12391
rect 20812 12238 20878 12391
rect 21004 12238 21070 12391
rect 21196 12238 21262 12391
rect 21388 12238 21454 12391
rect 21580 12238 21636 12391
rect 32 11737 98 11890
rect 224 11737 290 11890
rect 416 11737 482 11890
rect 608 11737 674 11890
rect 800 11737 866 11890
rect 992 11737 1058 11890
rect 1184 11737 1250 11890
rect 1376 11737 1442 11890
rect 1860 11737 1926 11890
rect 2052 11737 2118 11890
rect 2244 11737 2310 11890
rect 2436 11737 2502 11890
rect 2628 11737 2694 11890
rect 2820 11737 2886 11890
rect 3012 11737 3078 11890
rect 3204 11737 3270 11890
rect 3688 11737 3754 11890
rect 3880 11737 3946 11890
rect 4072 11737 4138 11890
rect 4264 11737 4330 11890
rect 4456 11737 4522 11890
rect 4648 11737 4714 11890
rect 4840 11737 4906 11890
rect 5032 11737 5098 11890
rect 5516 11737 5582 11890
rect 5708 11737 5774 11890
rect 5900 11737 5966 11890
rect 6092 11737 6158 11890
rect 6284 11737 6350 11890
rect 6476 11737 6542 11890
rect 6668 11737 6734 11890
rect 6860 11737 6926 11890
rect 7344 11737 7410 11890
rect 7536 11737 7602 11890
rect 7728 11737 7794 11890
rect 7920 11737 7986 11890
rect 8112 11737 8178 11890
rect 8304 11737 8370 11890
rect 8496 11737 8562 11890
rect 8688 11737 8754 11890
rect 9172 11737 9238 11890
rect 9364 11737 9430 11890
rect 9556 11737 9622 11890
rect 9748 11737 9814 11890
rect 9940 11737 10006 11890
rect 10132 11737 10198 11890
rect 10324 11737 10390 11890
rect 10516 11737 10582 11890
rect 11000 11737 11066 11890
rect 11192 11737 11258 11890
rect 11384 11737 11450 11890
rect 11576 11737 11642 11890
rect 11768 11737 11834 11890
rect 11960 11737 12026 11890
rect 12152 11737 12218 11890
rect 12344 11737 12410 11890
rect 12828 11737 12894 11890
rect 13020 11737 13086 11890
rect 13212 11737 13278 11890
rect 13404 11737 13470 11890
rect 13596 11737 13662 11890
rect 13788 11737 13854 11890
rect 13980 11737 14046 11890
rect 14172 11737 14238 11890
rect 14656 11737 14722 11890
rect 14848 11737 14914 11890
rect 15040 11737 15106 11890
rect 15232 11737 15298 11890
rect 15424 11737 15490 11890
rect 15616 11737 15682 11890
rect 15808 11737 15874 11890
rect 16000 11737 16066 11890
rect 16484 11737 16550 11890
rect 16676 11737 16742 11890
rect 16868 11737 16934 11890
rect 17060 11737 17126 11890
rect 17252 11737 17318 11890
rect 17444 11737 17510 11890
rect 17636 11737 17702 11890
rect 17828 11737 17894 11890
rect 18312 11737 18378 11890
rect 18504 11737 18570 11890
rect 18696 11737 18762 11890
rect 18888 11737 18954 11890
rect 19080 11737 19146 11890
rect 19272 11737 19338 11890
rect 19464 11737 19530 11890
rect 19656 11737 19722 11890
rect 20140 11737 20206 11890
rect 20332 11737 20398 11890
rect 20524 11737 20590 11890
rect 20716 11737 20782 11890
rect 20908 11737 20974 11890
rect 21100 11737 21166 11890
rect 21292 11737 21358 11890
rect 21484 11737 21550 11890
rect 128 11524 194 11677
rect 320 11524 386 11677
rect 512 11524 578 11677
rect 704 11524 770 11677
rect 896 11524 962 11677
rect 1088 11524 1154 11677
rect 1280 11524 1346 11677
rect 1472 11524 1528 11677
rect 1956 11524 2022 11677
rect 2148 11524 2214 11677
rect 2340 11524 2406 11677
rect 2532 11524 2598 11677
rect 2724 11524 2790 11677
rect 2916 11524 2982 11677
rect 3108 11524 3174 11677
rect 3300 11524 3356 11677
rect 3784 11524 3850 11677
rect 3976 11524 4042 11677
rect 4168 11524 4234 11677
rect 4360 11524 4426 11677
rect 4552 11524 4618 11677
rect 4744 11524 4810 11677
rect 4936 11524 5002 11677
rect 5128 11524 5184 11677
rect 5612 11524 5678 11677
rect 5804 11524 5870 11677
rect 5996 11524 6062 11677
rect 6188 11524 6254 11677
rect 6380 11524 6446 11677
rect 6572 11524 6638 11677
rect 6764 11524 6830 11677
rect 6956 11524 7012 11677
rect 7440 11524 7506 11677
rect 7632 11524 7698 11677
rect 7824 11524 7890 11677
rect 8016 11524 8082 11677
rect 8208 11524 8274 11677
rect 8400 11524 8466 11677
rect 8592 11524 8658 11677
rect 8784 11524 8840 11677
rect 9268 11524 9334 11677
rect 9460 11524 9526 11677
rect 9652 11524 9718 11677
rect 9844 11524 9910 11677
rect 10036 11524 10102 11677
rect 10228 11524 10294 11677
rect 10420 11524 10486 11677
rect 10612 11524 10668 11677
rect 11096 11524 11162 11677
rect 11288 11524 11354 11677
rect 11480 11524 11546 11677
rect 11672 11524 11738 11677
rect 11864 11524 11930 11677
rect 12056 11524 12122 11677
rect 12248 11524 12314 11677
rect 12440 11524 12496 11677
rect 12924 11524 12990 11677
rect 13116 11524 13182 11677
rect 13308 11524 13374 11677
rect 13500 11524 13566 11677
rect 13692 11524 13758 11677
rect 13884 11524 13950 11677
rect 14076 11524 14142 11677
rect 14268 11524 14324 11677
rect 14752 11524 14818 11677
rect 14944 11524 15010 11677
rect 15136 11524 15202 11677
rect 15328 11524 15394 11677
rect 15520 11524 15586 11677
rect 15712 11524 15778 11677
rect 15904 11524 15970 11677
rect 16096 11524 16152 11677
rect 16580 11524 16646 11677
rect 16772 11524 16838 11677
rect 16964 11524 17030 11677
rect 17156 11524 17222 11677
rect 17348 11524 17414 11677
rect 17540 11524 17606 11677
rect 17732 11524 17798 11677
rect 17924 11524 17980 11677
rect 18408 11524 18474 11677
rect 18600 11524 18666 11677
rect 18792 11524 18858 11677
rect 18984 11524 19050 11677
rect 19176 11524 19242 11677
rect 19368 11524 19434 11677
rect 19560 11524 19626 11677
rect 19752 11524 19808 11677
rect 20236 11524 20302 11677
rect 20428 11524 20494 11677
rect 20620 11524 20686 11677
rect 20812 11524 20878 11677
rect 21004 11524 21070 11677
rect 21196 11524 21262 11677
rect 21388 11524 21454 11677
rect 21580 11524 21636 11677
rect 32 11023 98 11176
rect 224 11023 290 11176
rect 416 11023 482 11176
rect 608 11023 674 11176
rect 800 11023 866 11176
rect 992 11023 1058 11176
rect 1184 11023 1250 11176
rect 1376 11023 1442 11176
rect 1860 11023 1926 11176
rect 2052 11023 2118 11176
rect 2244 11023 2310 11176
rect 2436 11023 2502 11176
rect 2628 11023 2694 11176
rect 2820 11023 2886 11176
rect 3012 11023 3078 11176
rect 3204 11023 3270 11176
rect 3688 11023 3754 11176
rect 3880 11023 3946 11176
rect 4072 11023 4138 11176
rect 4264 11023 4330 11176
rect 4456 11023 4522 11176
rect 4648 11023 4714 11176
rect 4840 11023 4906 11176
rect 5032 11023 5098 11176
rect 5516 11023 5582 11176
rect 5708 11023 5774 11176
rect 5900 11023 5966 11176
rect 6092 11023 6158 11176
rect 6284 11023 6350 11176
rect 6476 11023 6542 11176
rect 6668 11023 6734 11176
rect 6860 11023 6926 11176
rect 7344 11023 7410 11176
rect 7536 11023 7602 11176
rect 7728 11023 7794 11176
rect 7920 11023 7986 11176
rect 8112 11023 8178 11176
rect 8304 11023 8370 11176
rect 8496 11023 8562 11176
rect 8688 11023 8754 11176
rect 9172 11023 9238 11176
rect 9364 11023 9430 11176
rect 9556 11023 9622 11176
rect 9748 11023 9814 11176
rect 9940 11023 10006 11176
rect 10132 11023 10198 11176
rect 10324 11023 10390 11176
rect 10516 11023 10582 11176
rect 11000 11023 11066 11176
rect 11192 11023 11258 11176
rect 11384 11023 11450 11176
rect 11576 11023 11642 11176
rect 11768 11023 11834 11176
rect 11960 11023 12026 11176
rect 12152 11023 12218 11176
rect 12344 11023 12410 11176
rect 12828 11023 12894 11176
rect 13020 11023 13086 11176
rect 13212 11023 13278 11176
rect 13404 11023 13470 11176
rect 13596 11023 13662 11176
rect 13788 11023 13854 11176
rect 13980 11023 14046 11176
rect 14172 11023 14238 11176
rect 14656 11023 14722 11176
rect 14848 11023 14914 11176
rect 15040 11023 15106 11176
rect 15232 11023 15298 11176
rect 15424 11023 15490 11176
rect 15616 11023 15682 11176
rect 15808 11023 15874 11176
rect 16000 11023 16066 11176
rect 16484 11023 16550 11176
rect 16676 11023 16742 11176
rect 16868 11023 16934 11176
rect 17060 11023 17126 11176
rect 17252 11023 17318 11176
rect 17444 11023 17510 11176
rect 17636 11023 17702 11176
rect 17828 11023 17894 11176
rect 18312 11023 18378 11176
rect 18504 11023 18570 11176
rect 18696 11023 18762 11176
rect 18888 11023 18954 11176
rect 19080 11023 19146 11176
rect 19272 11023 19338 11176
rect 19464 11023 19530 11176
rect 19656 11023 19722 11176
rect 20140 11023 20206 11176
rect 20332 11023 20398 11176
rect 20524 11023 20590 11176
rect 20716 11023 20782 11176
rect 20908 11023 20974 11176
rect 21100 11023 21166 11176
rect 21292 11023 21358 11176
rect 21484 11023 21550 11176
rect 128 10810 194 10963
rect 320 10810 386 10963
rect 512 10810 578 10963
rect 704 10810 770 10963
rect 896 10810 962 10963
rect 1088 10810 1154 10963
rect 1280 10810 1346 10963
rect 1472 10810 1528 10963
rect 1956 10810 2022 10963
rect 2148 10810 2214 10963
rect 2340 10810 2406 10963
rect 2532 10810 2598 10963
rect 2724 10810 2790 10963
rect 2916 10810 2982 10963
rect 3108 10810 3174 10963
rect 3300 10810 3356 10963
rect 3784 10810 3850 10963
rect 3976 10810 4042 10963
rect 4168 10810 4234 10963
rect 4360 10810 4426 10963
rect 4552 10810 4618 10963
rect 4744 10810 4810 10963
rect 4936 10810 5002 10963
rect 5128 10810 5184 10963
rect 5612 10810 5678 10963
rect 5804 10810 5870 10963
rect 5996 10810 6062 10963
rect 6188 10810 6254 10963
rect 6380 10810 6446 10963
rect 6572 10810 6638 10963
rect 6764 10810 6830 10963
rect 6956 10810 7012 10963
rect 7440 10810 7506 10963
rect 7632 10810 7698 10963
rect 7824 10810 7890 10963
rect 8016 10810 8082 10963
rect 8208 10810 8274 10963
rect 8400 10810 8466 10963
rect 8592 10810 8658 10963
rect 8784 10810 8840 10963
rect 9268 10810 9334 10963
rect 9460 10810 9526 10963
rect 9652 10810 9718 10963
rect 9844 10810 9910 10963
rect 10036 10810 10102 10963
rect 10228 10810 10294 10963
rect 10420 10810 10486 10963
rect 10612 10810 10668 10963
rect 11096 10810 11162 10963
rect 11288 10810 11354 10963
rect 11480 10810 11546 10963
rect 11672 10810 11738 10963
rect 11864 10810 11930 10963
rect 12056 10810 12122 10963
rect 12248 10810 12314 10963
rect 12440 10810 12496 10963
rect 12924 10810 12990 10963
rect 13116 10810 13182 10963
rect 13308 10810 13374 10963
rect 13500 10810 13566 10963
rect 13692 10810 13758 10963
rect 13884 10810 13950 10963
rect 14076 10810 14142 10963
rect 14268 10810 14324 10963
rect 14752 10810 14818 10963
rect 14944 10810 15010 10963
rect 15136 10810 15202 10963
rect 15328 10810 15394 10963
rect 15520 10810 15586 10963
rect 15712 10810 15778 10963
rect 15904 10810 15970 10963
rect 16096 10810 16152 10963
rect 16580 10810 16646 10963
rect 16772 10810 16838 10963
rect 16964 10810 17030 10963
rect 17156 10810 17222 10963
rect 17348 10810 17414 10963
rect 17540 10810 17606 10963
rect 17732 10810 17798 10963
rect 17924 10810 17980 10963
rect 18408 10810 18474 10963
rect 18600 10810 18666 10963
rect 18792 10810 18858 10963
rect 18984 10810 19050 10963
rect 19176 10810 19242 10963
rect 19368 10810 19434 10963
rect 19560 10810 19626 10963
rect 19752 10810 19808 10963
rect 20236 10810 20302 10963
rect 20428 10810 20494 10963
rect 20620 10810 20686 10963
rect 20812 10810 20878 10963
rect 21004 10810 21070 10963
rect 21196 10810 21262 10963
rect 21388 10810 21454 10963
rect 21580 10810 21636 10963
rect 32 10309 98 10462
rect 224 10309 290 10462
rect 416 10309 482 10462
rect 608 10309 674 10462
rect 800 10309 866 10462
rect 992 10309 1058 10462
rect 1184 10309 1250 10462
rect 1376 10309 1442 10462
rect 1860 10309 1926 10462
rect 2052 10309 2118 10462
rect 2244 10309 2310 10462
rect 2436 10309 2502 10462
rect 2628 10309 2694 10462
rect 2820 10309 2886 10462
rect 3012 10309 3078 10462
rect 3204 10309 3270 10462
rect 3688 10309 3754 10462
rect 3880 10309 3946 10462
rect 4072 10309 4138 10462
rect 4264 10309 4330 10462
rect 4456 10309 4522 10462
rect 4648 10309 4714 10462
rect 4840 10309 4906 10462
rect 5032 10309 5098 10462
rect 5516 10309 5582 10462
rect 5708 10309 5774 10462
rect 5900 10309 5966 10462
rect 6092 10309 6158 10462
rect 6284 10309 6350 10462
rect 6476 10309 6542 10462
rect 6668 10309 6734 10462
rect 6860 10309 6926 10462
rect 7344 10309 7410 10462
rect 7536 10309 7602 10462
rect 7728 10309 7794 10462
rect 7920 10309 7986 10462
rect 8112 10309 8178 10462
rect 8304 10309 8370 10462
rect 8496 10309 8562 10462
rect 8688 10309 8754 10462
rect 9172 10309 9238 10462
rect 9364 10309 9430 10462
rect 9556 10309 9622 10462
rect 9748 10309 9814 10462
rect 9940 10309 10006 10462
rect 10132 10309 10198 10462
rect 10324 10309 10390 10462
rect 10516 10309 10582 10462
rect 11000 10309 11066 10462
rect 11192 10309 11258 10462
rect 11384 10309 11450 10462
rect 11576 10309 11642 10462
rect 11768 10309 11834 10462
rect 11960 10309 12026 10462
rect 12152 10309 12218 10462
rect 12344 10309 12410 10462
rect 12828 10309 12894 10462
rect 13020 10309 13086 10462
rect 13212 10309 13278 10462
rect 13404 10309 13470 10462
rect 13596 10309 13662 10462
rect 13788 10309 13854 10462
rect 13980 10309 14046 10462
rect 14172 10309 14238 10462
rect 14656 10309 14722 10462
rect 14848 10309 14914 10462
rect 15040 10309 15106 10462
rect 15232 10309 15298 10462
rect 15424 10309 15490 10462
rect 15616 10309 15682 10462
rect 15808 10309 15874 10462
rect 16000 10309 16066 10462
rect 16484 10309 16550 10462
rect 16676 10309 16742 10462
rect 16868 10309 16934 10462
rect 17060 10309 17126 10462
rect 17252 10309 17318 10462
rect 17444 10309 17510 10462
rect 17636 10309 17702 10462
rect 17828 10309 17894 10462
rect 18312 10309 18378 10462
rect 18504 10309 18570 10462
rect 18696 10309 18762 10462
rect 18888 10309 18954 10462
rect 19080 10309 19146 10462
rect 19272 10309 19338 10462
rect 19464 10309 19530 10462
rect 19656 10309 19722 10462
rect 20140 10309 20206 10462
rect 20332 10309 20398 10462
rect 20524 10309 20590 10462
rect 20716 10309 20782 10462
rect 20908 10309 20974 10462
rect 21100 10309 21166 10462
rect 21292 10309 21358 10462
rect 21484 10309 21550 10462
rect 128 10096 194 10249
rect 320 10096 386 10249
rect 512 10096 578 10249
rect 704 10096 770 10249
rect 896 10096 962 10249
rect 1088 10096 1154 10249
rect 1280 10096 1346 10249
rect 1472 10096 1528 10249
rect 1956 10096 2022 10249
rect 2148 10096 2214 10249
rect 2340 10096 2406 10249
rect 2532 10096 2598 10249
rect 2724 10096 2790 10249
rect 2916 10096 2982 10249
rect 3108 10096 3174 10249
rect 3300 10096 3356 10249
rect 3784 10096 3850 10249
rect 3976 10096 4042 10249
rect 4168 10096 4234 10249
rect 4360 10096 4426 10249
rect 4552 10096 4618 10249
rect 4744 10096 4810 10249
rect 4936 10096 5002 10249
rect 5128 10096 5184 10249
rect 5612 10096 5678 10249
rect 5804 10096 5870 10249
rect 5996 10096 6062 10249
rect 6188 10096 6254 10249
rect 6380 10096 6446 10249
rect 6572 10096 6638 10249
rect 6764 10096 6830 10249
rect 6956 10096 7012 10249
rect 7440 10096 7506 10249
rect 7632 10096 7698 10249
rect 7824 10096 7890 10249
rect 8016 10096 8082 10249
rect 8208 10096 8274 10249
rect 8400 10096 8466 10249
rect 8592 10096 8658 10249
rect 8784 10096 8840 10249
rect 9268 10096 9334 10249
rect 9460 10096 9526 10249
rect 9652 10096 9718 10249
rect 9844 10096 9910 10249
rect 10036 10096 10102 10249
rect 10228 10096 10294 10249
rect 10420 10096 10486 10249
rect 10612 10096 10668 10249
rect 11096 10096 11162 10249
rect 11288 10096 11354 10249
rect 11480 10096 11546 10249
rect 11672 10096 11738 10249
rect 11864 10096 11930 10249
rect 12056 10096 12122 10249
rect 12248 10096 12314 10249
rect 12440 10096 12496 10249
rect 12924 10096 12990 10249
rect 13116 10096 13182 10249
rect 13308 10096 13374 10249
rect 13500 10096 13566 10249
rect 13692 10096 13758 10249
rect 13884 10096 13950 10249
rect 14076 10096 14142 10249
rect 14268 10096 14324 10249
rect 14752 10096 14818 10249
rect 14944 10096 15010 10249
rect 15136 10096 15202 10249
rect 15328 10096 15394 10249
rect 15520 10096 15586 10249
rect 15712 10096 15778 10249
rect 15904 10096 15970 10249
rect 16096 10096 16152 10249
rect 16580 10096 16646 10249
rect 16772 10096 16838 10249
rect 16964 10096 17030 10249
rect 17156 10096 17222 10249
rect 17348 10096 17414 10249
rect 17540 10096 17606 10249
rect 17732 10096 17798 10249
rect 17924 10096 17980 10249
rect 18408 10096 18474 10249
rect 18600 10096 18666 10249
rect 18792 10096 18858 10249
rect 18984 10096 19050 10249
rect 19176 10096 19242 10249
rect 19368 10096 19434 10249
rect 19560 10096 19626 10249
rect 19752 10096 19808 10249
rect 20236 10096 20302 10249
rect 20428 10096 20494 10249
rect 20620 10096 20686 10249
rect 20812 10096 20878 10249
rect 21004 10096 21070 10249
rect 21196 10096 21262 10249
rect 21388 10096 21454 10249
rect 21580 10096 21636 10249
rect 32 9595 98 9748
rect 224 9595 290 9748
rect 416 9595 482 9748
rect 608 9595 674 9748
rect 800 9595 866 9748
rect 992 9595 1058 9748
rect 1184 9595 1250 9748
rect 1376 9595 1442 9748
rect 1860 9595 1926 9748
rect 2052 9595 2118 9748
rect 2244 9595 2310 9748
rect 2436 9595 2502 9748
rect 2628 9595 2694 9748
rect 2820 9595 2886 9748
rect 3012 9595 3078 9748
rect 3204 9595 3270 9748
rect 3688 9595 3754 9748
rect 3880 9595 3946 9748
rect 4072 9595 4138 9748
rect 4264 9595 4330 9748
rect 4456 9595 4522 9748
rect 4648 9595 4714 9748
rect 4840 9595 4906 9748
rect 5032 9595 5098 9748
rect 5516 9595 5582 9748
rect 5708 9595 5774 9748
rect 5900 9595 5966 9748
rect 6092 9595 6158 9748
rect 6284 9595 6350 9748
rect 6476 9595 6542 9748
rect 6668 9595 6734 9748
rect 6860 9595 6926 9748
rect 7344 9595 7410 9748
rect 7536 9595 7602 9748
rect 7728 9595 7794 9748
rect 7920 9595 7986 9748
rect 8112 9595 8178 9748
rect 8304 9595 8370 9748
rect 8496 9595 8562 9748
rect 8688 9595 8754 9748
rect 9172 9595 9238 9748
rect 9364 9595 9430 9748
rect 9556 9595 9622 9748
rect 9748 9595 9814 9748
rect 9940 9595 10006 9748
rect 10132 9595 10198 9748
rect 10324 9595 10390 9748
rect 10516 9595 10582 9748
rect 11000 9595 11066 9748
rect 11192 9595 11258 9748
rect 11384 9595 11450 9748
rect 11576 9595 11642 9748
rect 11768 9595 11834 9748
rect 11960 9595 12026 9748
rect 12152 9595 12218 9748
rect 12344 9595 12410 9748
rect 12828 9595 12894 9748
rect 13020 9595 13086 9748
rect 13212 9595 13278 9748
rect 13404 9595 13470 9748
rect 13596 9595 13662 9748
rect 13788 9595 13854 9748
rect 13980 9595 14046 9748
rect 14172 9595 14238 9748
rect 14656 9595 14722 9748
rect 14848 9595 14914 9748
rect 15040 9595 15106 9748
rect 15232 9595 15298 9748
rect 15424 9595 15490 9748
rect 15616 9595 15682 9748
rect 15808 9595 15874 9748
rect 16000 9595 16066 9748
rect 16484 9595 16550 9748
rect 16676 9595 16742 9748
rect 16868 9595 16934 9748
rect 17060 9595 17126 9748
rect 17252 9595 17318 9748
rect 17444 9595 17510 9748
rect 17636 9595 17702 9748
rect 17828 9595 17894 9748
rect 18312 9595 18378 9748
rect 18504 9595 18570 9748
rect 18696 9595 18762 9748
rect 18888 9595 18954 9748
rect 19080 9595 19146 9748
rect 19272 9595 19338 9748
rect 19464 9595 19530 9748
rect 19656 9595 19722 9748
rect 20140 9595 20206 9748
rect 20332 9595 20398 9748
rect 20524 9595 20590 9748
rect 20716 9595 20782 9748
rect 20908 9595 20974 9748
rect 21100 9595 21166 9748
rect 21292 9595 21358 9748
rect 21484 9595 21550 9748
rect 128 9382 194 9535
rect 320 9382 386 9535
rect 512 9382 578 9535
rect 704 9382 770 9535
rect 896 9382 962 9535
rect 1088 9382 1154 9535
rect 1280 9382 1346 9535
rect 1472 9382 1528 9535
rect 1956 9382 2022 9535
rect 2148 9382 2214 9535
rect 2340 9382 2406 9535
rect 2532 9382 2598 9535
rect 2724 9382 2790 9535
rect 2916 9382 2982 9535
rect 3108 9382 3174 9535
rect 3300 9382 3356 9535
rect 3784 9382 3850 9535
rect 3976 9382 4042 9535
rect 4168 9382 4234 9535
rect 4360 9382 4426 9535
rect 4552 9382 4618 9535
rect 4744 9382 4810 9535
rect 4936 9382 5002 9535
rect 5128 9382 5184 9535
rect 5612 9382 5678 9535
rect 5804 9382 5870 9535
rect 5996 9382 6062 9535
rect 6188 9382 6254 9535
rect 6380 9382 6446 9535
rect 6572 9382 6638 9535
rect 6764 9382 6830 9535
rect 6956 9382 7012 9535
rect 7440 9382 7506 9535
rect 7632 9382 7698 9535
rect 7824 9382 7890 9535
rect 8016 9382 8082 9535
rect 8208 9382 8274 9535
rect 8400 9382 8466 9535
rect 8592 9382 8658 9535
rect 8784 9382 8840 9535
rect 9268 9382 9334 9535
rect 9460 9382 9526 9535
rect 9652 9382 9718 9535
rect 9844 9382 9910 9535
rect 10036 9382 10102 9535
rect 10228 9382 10294 9535
rect 10420 9382 10486 9535
rect 10612 9382 10668 9535
rect 11096 9382 11162 9535
rect 11288 9382 11354 9535
rect 11480 9382 11546 9535
rect 11672 9382 11738 9535
rect 11864 9382 11930 9535
rect 12056 9382 12122 9535
rect 12248 9382 12314 9535
rect 12440 9382 12496 9535
rect 12924 9382 12990 9535
rect 13116 9382 13182 9535
rect 13308 9382 13374 9535
rect 13500 9382 13566 9535
rect 13692 9382 13758 9535
rect 13884 9382 13950 9535
rect 14076 9382 14142 9535
rect 14268 9382 14324 9535
rect 14752 9382 14818 9535
rect 14944 9382 15010 9535
rect 15136 9382 15202 9535
rect 15328 9382 15394 9535
rect 15520 9382 15586 9535
rect 15712 9382 15778 9535
rect 15904 9382 15970 9535
rect 16096 9382 16152 9535
rect 16580 9382 16646 9535
rect 16772 9382 16838 9535
rect 16964 9382 17030 9535
rect 17156 9382 17222 9535
rect 17348 9382 17414 9535
rect 17540 9382 17606 9535
rect 17732 9382 17798 9535
rect 17924 9382 17980 9535
rect 18408 9382 18474 9535
rect 18600 9382 18666 9535
rect 18792 9382 18858 9535
rect 18984 9382 19050 9535
rect 19176 9382 19242 9535
rect 19368 9382 19434 9535
rect 19560 9382 19626 9535
rect 19752 9382 19808 9535
rect 20236 9382 20302 9535
rect 20428 9382 20494 9535
rect 20620 9382 20686 9535
rect 20812 9382 20878 9535
rect 21004 9382 21070 9535
rect 21196 9382 21262 9535
rect 21388 9382 21454 9535
rect 21580 9382 21636 9535
rect 32 8881 98 9034
rect 224 8881 290 9034
rect 416 8881 482 9034
rect 608 8881 674 9034
rect 800 8881 866 9034
rect 992 8881 1058 9034
rect 1184 8881 1250 9034
rect 1376 8881 1442 9034
rect 1860 8881 1926 9034
rect 2052 8881 2118 9034
rect 2244 8881 2310 9034
rect 2436 8881 2502 9034
rect 2628 8881 2694 9034
rect 2820 8881 2886 9034
rect 3012 8881 3078 9034
rect 3204 8881 3270 9034
rect 3688 8881 3754 9034
rect 3880 8881 3946 9034
rect 4072 8881 4138 9034
rect 4264 8881 4330 9034
rect 4456 8881 4522 9034
rect 4648 8881 4714 9034
rect 4840 8881 4906 9034
rect 5032 8881 5098 9034
rect 5516 8881 5582 9034
rect 5708 8881 5774 9034
rect 5900 8881 5966 9034
rect 6092 8881 6158 9034
rect 6284 8881 6350 9034
rect 6476 8881 6542 9034
rect 6668 8881 6734 9034
rect 6860 8881 6926 9034
rect 7344 8881 7410 9034
rect 7536 8881 7602 9034
rect 7728 8881 7794 9034
rect 7920 8881 7986 9034
rect 8112 8881 8178 9034
rect 8304 8881 8370 9034
rect 8496 8881 8562 9034
rect 8688 8881 8754 9034
rect 9172 8881 9238 9034
rect 9364 8881 9430 9034
rect 9556 8881 9622 9034
rect 9748 8881 9814 9034
rect 9940 8881 10006 9034
rect 10132 8881 10198 9034
rect 10324 8881 10390 9034
rect 10516 8881 10582 9034
rect 11000 8881 11066 9034
rect 11192 8881 11258 9034
rect 11384 8881 11450 9034
rect 11576 8881 11642 9034
rect 11768 8881 11834 9034
rect 11960 8881 12026 9034
rect 12152 8881 12218 9034
rect 12344 8881 12410 9034
rect 12828 8881 12894 9034
rect 13020 8881 13086 9034
rect 13212 8881 13278 9034
rect 13404 8881 13470 9034
rect 13596 8881 13662 9034
rect 13788 8881 13854 9034
rect 13980 8881 14046 9034
rect 14172 8881 14238 9034
rect 14656 8881 14722 9034
rect 14848 8881 14914 9034
rect 15040 8881 15106 9034
rect 15232 8881 15298 9034
rect 15424 8881 15490 9034
rect 15616 8881 15682 9034
rect 15808 8881 15874 9034
rect 16000 8881 16066 9034
rect 16484 8881 16550 9034
rect 16676 8881 16742 9034
rect 16868 8881 16934 9034
rect 17060 8881 17126 9034
rect 17252 8881 17318 9034
rect 17444 8881 17510 9034
rect 17636 8881 17702 9034
rect 17828 8881 17894 9034
rect 18312 8881 18378 9034
rect 18504 8881 18570 9034
rect 18696 8881 18762 9034
rect 18888 8881 18954 9034
rect 19080 8881 19146 9034
rect 19272 8881 19338 9034
rect 19464 8881 19530 9034
rect 19656 8881 19722 9034
rect 20140 8881 20206 9034
rect 20332 8881 20398 9034
rect 20524 8881 20590 9034
rect 20716 8881 20782 9034
rect 20908 8881 20974 9034
rect 21100 8881 21166 9034
rect 21292 8881 21358 9034
rect 21484 8881 21550 9034
rect 128 8668 194 8821
rect 320 8668 386 8821
rect 512 8668 578 8821
rect 704 8668 770 8821
rect 896 8668 962 8821
rect 1088 8668 1154 8821
rect 1280 8668 1346 8821
rect 1472 8668 1528 8821
rect 1956 8668 2022 8821
rect 2148 8668 2214 8821
rect 2340 8668 2406 8821
rect 2532 8668 2598 8821
rect 2724 8668 2790 8821
rect 2916 8668 2982 8821
rect 3108 8668 3174 8821
rect 3300 8668 3356 8821
rect 3784 8668 3850 8821
rect 3976 8668 4042 8821
rect 4168 8668 4234 8821
rect 4360 8668 4426 8821
rect 4552 8668 4618 8821
rect 4744 8668 4810 8821
rect 4936 8668 5002 8821
rect 5128 8668 5184 8821
rect 5612 8668 5678 8821
rect 5804 8668 5870 8821
rect 5996 8668 6062 8821
rect 6188 8668 6254 8821
rect 6380 8668 6446 8821
rect 6572 8668 6638 8821
rect 6764 8668 6830 8821
rect 6956 8668 7012 8821
rect 7440 8668 7506 8821
rect 7632 8668 7698 8821
rect 7824 8668 7890 8821
rect 8016 8668 8082 8821
rect 8208 8668 8274 8821
rect 8400 8668 8466 8821
rect 8592 8668 8658 8821
rect 8784 8668 8840 8821
rect 9268 8668 9334 8821
rect 9460 8668 9526 8821
rect 9652 8668 9718 8821
rect 9844 8668 9910 8821
rect 10036 8668 10102 8821
rect 10228 8668 10294 8821
rect 10420 8668 10486 8821
rect 10612 8668 10668 8821
rect 11096 8668 11162 8821
rect 11288 8668 11354 8821
rect 11480 8668 11546 8821
rect 11672 8668 11738 8821
rect 11864 8668 11930 8821
rect 12056 8668 12122 8821
rect 12248 8668 12314 8821
rect 12440 8668 12496 8821
rect 12924 8668 12990 8821
rect 13116 8668 13182 8821
rect 13308 8668 13374 8821
rect 13500 8668 13566 8821
rect 13692 8668 13758 8821
rect 13884 8668 13950 8821
rect 14076 8668 14142 8821
rect 14268 8668 14324 8821
rect 14752 8668 14818 8821
rect 14944 8668 15010 8821
rect 15136 8668 15202 8821
rect 15328 8668 15394 8821
rect 15520 8668 15586 8821
rect 15712 8668 15778 8821
rect 15904 8668 15970 8821
rect 16096 8668 16152 8821
rect 16580 8668 16646 8821
rect 16772 8668 16838 8821
rect 16964 8668 17030 8821
rect 17156 8668 17222 8821
rect 17348 8668 17414 8821
rect 17540 8668 17606 8821
rect 17732 8668 17798 8821
rect 17924 8668 17980 8821
rect 18408 8668 18474 8821
rect 18600 8668 18666 8821
rect 18792 8668 18858 8821
rect 18984 8668 19050 8821
rect 19176 8668 19242 8821
rect 19368 8668 19434 8821
rect 19560 8668 19626 8821
rect 19752 8668 19808 8821
rect 20236 8668 20302 8821
rect 20428 8668 20494 8821
rect 20620 8668 20686 8821
rect 20812 8668 20878 8821
rect 21004 8668 21070 8821
rect 21196 8668 21262 8821
rect 21388 8668 21454 8821
rect 21580 8668 21636 8821
rect 32 8167 98 8320
rect 224 8167 290 8320
rect 416 8167 482 8320
rect 608 8167 674 8320
rect 800 8167 866 8320
rect 992 8167 1058 8320
rect 1184 8167 1250 8320
rect 1376 8167 1442 8320
rect 1860 8167 1926 8320
rect 2052 8167 2118 8320
rect 2244 8167 2310 8320
rect 2436 8167 2502 8320
rect 2628 8167 2694 8320
rect 2820 8167 2886 8320
rect 3012 8167 3078 8320
rect 3204 8167 3270 8320
rect 3688 8167 3754 8320
rect 3880 8167 3946 8320
rect 4072 8167 4138 8320
rect 4264 8167 4330 8320
rect 4456 8167 4522 8320
rect 4648 8167 4714 8320
rect 4840 8167 4906 8320
rect 5032 8167 5098 8320
rect 5516 8167 5582 8320
rect 5708 8167 5774 8320
rect 5900 8167 5966 8320
rect 6092 8167 6158 8320
rect 6284 8167 6350 8320
rect 6476 8167 6542 8320
rect 6668 8167 6734 8320
rect 6860 8167 6926 8320
rect 7344 8167 7410 8320
rect 7536 8167 7602 8320
rect 7728 8167 7794 8320
rect 7920 8167 7986 8320
rect 8112 8167 8178 8320
rect 8304 8167 8370 8320
rect 8496 8167 8562 8320
rect 8688 8167 8754 8320
rect 9172 8167 9238 8320
rect 9364 8167 9430 8320
rect 9556 8167 9622 8320
rect 9748 8167 9814 8320
rect 9940 8167 10006 8320
rect 10132 8167 10198 8320
rect 10324 8167 10390 8320
rect 10516 8167 10582 8320
rect 11000 8167 11066 8320
rect 11192 8167 11258 8320
rect 11384 8167 11450 8320
rect 11576 8167 11642 8320
rect 11768 8167 11834 8320
rect 11960 8167 12026 8320
rect 12152 8167 12218 8320
rect 12344 8167 12410 8320
rect 12828 8167 12894 8320
rect 13020 8167 13086 8320
rect 13212 8167 13278 8320
rect 13404 8167 13470 8320
rect 13596 8167 13662 8320
rect 13788 8167 13854 8320
rect 13980 8167 14046 8320
rect 14172 8167 14238 8320
rect 14656 8167 14722 8320
rect 14848 8167 14914 8320
rect 15040 8167 15106 8320
rect 15232 8167 15298 8320
rect 15424 8167 15490 8320
rect 15616 8167 15682 8320
rect 15808 8167 15874 8320
rect 16000 8167 16066 8320
rect 16484 8167 16550 8320
rect 16676 8167 16742 8320
rect 16868 8167 16934 8320
rect 17060 8167 17126 8320
rect 17252 8167 17318 8320
rect 17444 8167 17510 8320
rect 17636 8167 17702 8320
rect 17828 8167 17894 8320
rect 18312 8167 18378 8320
rect 18504 8167 18570 8320
rect 18696 8167 18762 8320
rect 18888 8167 18954 8320
rect 19080 8167 19146 8320
rect 19272 8167 19338 8320
rect 19464 8167 19530 8320
rect 19656 8167 19722 8320
rect 20140 8167 20206 8320
rect 20332 8167 20398 8320
rect 20524 8167 20590 8320
rect 20716 8167 20782 8320
rect 20908 8167 20974 8320
rect 21100 8167 21166 8320
rect 21292 8167 21358 8320
rect 21484 8167 21550 8320
rect 128 7954 194 8107
rect 320 7954 386 8107
rect 512 7954 578 8107
rect 704 7954 770 8107
rect 896 7954 962 8107
rect 1088 7954 1154 8107
rect 1280 7954 1346 8107
rect 1472 7954 1528 8107
rect 1956 7954 2022 8107
rect 2148 7954 2214 8107
rect 2340 7954 2406 8107
rect 2532 7954 2598 8107
rect 2724 7954 2790 8107
rect 2916 7954 2982 8107
rect 3108 7954 3174 8107
rect 3300 7954 3356 8107
rect 3784 7954 3850 8107
rect 3976 7954 4042 8107
rect 4168 7954 4234 8107
rect 4360 7954 4426 8107
rect 4552 7954 4618 8107
rect 4744 7954 4810 8107
rect 4936 7954 5002 8107
rect 5128 7954 5184 8107
rect 5612 7954 5678 8107
rect 5804 7954 5870 8107
rect 5996 7954 6062 8107
rect 6188 7954 6254 8107
rect 6380 7954 6446 8107
rect 6572 7954 6638 8107
rect 6764 7954 6830 8107
rect 6956 7954 7012 8107
rect 7440 7954 7506 8107
rect 7632 7954 7698 8107
rect 7824 7954 7890 8107
rect 8016 7954 8082 8107
rect 8208 7954 8274 8107
rect 8400 7954 8466 8107
rect 8592 7954 8658 8107
rect 8784 7954 8840 8107
rect 9268 7954 9334 8107
rect 9460 7954 9526 8107
rect 9652 7954 9718 8107
rect 9844 7954 9910 8107
rect 10036 7954 10102 8107
rect 10228 7954 10294 8107
rect 10420 7954 10486 8107
rect 10612 7954 10668 8107
rect 11096 7954 11162 8107
rect 11288 7954 11354 8107
rect 11480 7954 11546 8107
rect 11672 7954 11738 8107
rect 11864 7954 11930 8107
rect 12056 7954 12122 8107
rect 12248 7954 12314 8107
rect 12440 7954 12496 8107
rect 12924 7954 12990 8107
rect 13116 7954 13182 8107
rect 13308 7954 13374 8107
rect 13500 7954 13566 8107
rect 13692 7954 13758 8107
rect 13884 7954 13950 8107
rect 14076 7954 14142 8107
rect 14268 7954 14324 8107
rect 14752 7954 14818 8107
rect 14944 7954 15010 8107
rect 15136 7954 15202 8107
rect 15328 7954 15394 8107
rect 15520 7954 15586 8107
rect 15712 7954 15778 8107
rect 15904 7954 15970 8107
rect 16096 7954 16152 8107
rect 16580 7954 16646 8107
rect 16772 7954 16838 8107
rect 16964 7954 17030 8107
rect 17156 7954 17222 8107
rect 17348 7954 17414 8107
rect 17540 7954 17606 8107
rect 17732 7954 17798 8107
rect 17924 7954 17980 8107
rect 18408 7954 18474 8107
rect 18600 7954 18666 8107
rect 18792 7954 18858 8107
rect 18984 7954 19050 8107
rect 19176 7954 19242 8107
rect 19368 7954 19434 8107
rect 19560 7954 19626 8107
rect 19752 7954 19808 8107
rect 20236 7954 20302 8107
rect 20428 7954 20494 8107
rect 20620 7954 20686 8107
rect 20812 7954 20878 8107
rect 21004 7954 21070 8107
rect 21196 7954 21262 8107
rect 21388 7954 21454 8107
rect 21580 7954 21636 8107
rect 32 7453 98 7606
rect 224 7453 290 7606
rect 416 7453 482 7606
rect 608 7453 674 7606
rect 800 7453 866 7606
rect 992 7453 1058 7606
rect 1184 7453 1250 7606
rect 1376 7453 1442 7606
rect 1860 7453 1926 7606
rect 2052 7453 2118 7606
rect 2244 7453 2310 7606
rect 2436 7453 2502 7606
rect 2628 7453 2694 7606
rect 2820 7453 2886 7606
rect 3012 7453 3078 7606
rect 3204 7453 3270 7606
rect 3688 7453 3754 7606
rect 3880 7453 3946 7606
rect 4072 7453 4138 7606
rect 4264 7453 4330 7606
rect 4456 7453 4522 7606
rect 4648 7453 4714 7606
rect 4840 7453 4906 7606
rect 5032 7453 5098 7606
rect 5516 7453 5582 7606
rect 5708 7453 5774 7606
rect 5900 7453 5966 7606
rect 6092 7453 6158 7606
rect 6284 7453 6350 7606
rect 6476 7453 6542 7606
rect 6668 7453 6734 7606
rect 6860 7453 6926 7606
rect 7344 7453 7410 7606
rect 7536 7453 7602 7606
rect 7728 7453 7794 7606
rect 7920 7453 7986 7606
rect 8112 7453 8178 7606
rect 8304 7453 8370 7606
rect 8496 7453 8562 7606
rect 8688 7453 8754 7606
rect 9172 7453 9238 7606
rect 9364 7453 9430 7606
rect 9556 7453 9622 7606
rect 9748 7453 9814 7606
rect 9940 7453 10006 7606
rect 10132 7453 10198 7606
rect 10324 7453 10390 7606
rect 10516 7453 10582 7606
rect 11000 7453 11066 7606
rect 11192 7453 11258 7606
rect 11384 7453 11450 7606
rect 11576 7453 11642 7606
rect 11768 7453 11834 7606
rect 11960 7453 12026 7606
rect 12152 7453 12218 7606
rect 12344 7453 12410 7606
rect 12828 7453 12894 7606
rect 13020 7453 13086 7606
rect 13212 7453 13278 7606
rect 13404 7453 13470 7606
rect 13596 7453 13662 7606
rect 13788 7453 13854 7606
rect 13980 7453 14046 7606
rect 14172 7453 14238 7606
rect 14656 7453 14722 7606
rect 14848 7453 14914 7606
rect 15040 7453 15106 7606
rect 15232 7453 15298 7606
rect 15424 7453 15490 7606
rect 15616 7453 15682 7606
rect 15808 7453 15874 7606
rect 16000 7453 16066 7606
rect 16484 7453 16550 7606
rect 16676 7453 16742 7606
rect 16868 7453 16934 7606
rect 17060 7453 17126 7606
rect 17252 7453 17318 7606
rect 17444 7453 17510 7606
rect 17636 7453 17702 7606
rect 17828 7453 17894 7606
rect 18312 7453 18378 7606
rect 18504 7453 18570 7606
rect 18696 7453 18762 7606
rect 18888 7453 18954 7606
rect 19080 7453 19146 7606
rect 19272 7453 19338 7606
rect 19464 7453 19530 7606
rect 19656 7453 19722 7606
rect 20140 7453 20206 7606
rect 20332 7453 20398 7606
rect 20524 7453 20590 7606
rect 20716 7453 20782 7606
rect 20908 7453 20974 7606
rect 21100 7453 21166 7606
rect 21292 7453 21358 7606
rect 21484 7453 21550 7606
rect 128 7240 194 7393
rect 320 7240 386 7393
rect 512 7240 578 7393
rect 704 7240 770 7393
rect 896 7240 962 7393
rect 1088 7240 1154 7393
rect 1280 7240 1346 7393
rect 1472 7240 1528 7393
rect 1956 7240 2022 7393
rect 2148 7240 2214 7393
rect 2340 7240 2406 7393
rect 2532 7240 2598 7393
rect 2724 7240 2790 7393
rect 2916 7240 2982 7393
rect 3108 7240 3174 7393
rect 3300 7240 3356 7393
rect 3784 7240 3850 7393
rect 3976 7240 4042 7393
rect 4168 7240 4234 7393
rect 4360 7240 4426 7393
rect 4552 7240 4618 7393
rect 4744 7240 4810 7393
rect 4936 7240 5002 7393
rect 5128 7240 5184 7393
rect 5612 7240 5678 7393
rect 5804 7240 5870 7393
rect 5996 7240 6062 7393
rect 6188 7240 6254 7393
rect 6380 7240 6446 7393
rect 6572 7240 6638 7393
rect 6764 7240 6830 7393
rect 6956 7240 7012 7393
rect 7440 7240 7506 7393
rect 7632 7240 7698 7393
rect 7824 7240 7890 7393
rect 8016 7240 8082 7393
rect 8208 7240 8274 7393
rect 8400 7240 8466 7393
rect 8592 7240 8658 7393
rect 8784 7240 8840 7393
rect 9268 7240 9334 7393
rect 9460 7240 9526 7393
rect 9652 7240 9718 7393
rect 9844 7240 9910 7393
rect 10036 7240 10102 7393
rect 10228 7240 10294 7393
rect 10420 7240 10486 7393
rect 10612 7240 10668 7393
rect 11096 7240 11162 7393
rect 11288 7240 11354 7393
rect 11480 7240 11546 7393
rect 11672 7240 11738 7393
rect 11864 7240 11930 7393
rect 12056 7240 12122 7393
rect 12248 7240 12314 7393
rect 12440 7240 12496 7393
rect 12924 7240 12990 7393
rect 13116 7240 13182 7393
rect 13308 7240 13374 7393
rect 13500 7240 13566 7393
rect 13692 7240 13758 7393
rect 13884 7240 13950 7393
rect 14076 7240 14142 7393
rect 14268 7240 14324 7393
rect 14752 7240 14818 7393
rect 14944 7240 15010 7393
rect 15136 7240 15202 7393
rect 15328 7240 15394 7393
rect 15520 7240 15586 7393
rect 15712 7240 15778 7393
rect 15904 7240 15970 7393
rect 16096 7240 16152 7393
rect 16580 7240 16646 7393
rect 16772 7240 16838 7393
rect 16964 7240 17030 7393
rect 17156 7240 17222 7393
rect 17348 7240 17414 7393
rect 17540 7240 17606 7393
rect 17732 7240 17798 7393
rect 17924 7240 17980 7393
rect 18408 7240 18474 7393
rect 18600 7240 18666 7393
rect 18792 7240 18858 7393
rect 18984 7240 19050 7393
rect 19176 7240 19242 7393
rect 19368 7240 19434 7393
rect 19560 7240 19626 7393
rect 19752 7240 19808 7393
rect 20236 7240 20302 7393
rect 20428 7240 20494 7393
rect 20620 7240 20686 7393
rect 20812 7240 20878 7393
rect 21004 7240 21070 7393
rect 21196 7240 21262 7393
rect 21388 7240 21454 7393
rect 21580 7240 21636 7393
rect 32 6739 98 6892
rect 224 6739 290 6892
rect 416 6739 482 6892
rect 608 6739 674 6892
rect 800 6739 866 6892
rect 992 6739 1058 6892
rect 1184 6739 1250 6892
rect 1376 6739 1442 6892
rect 1860 6739 1926 6892
rect 2052 6739 2118 6892
rect 2244 6739 2310 6892
rect 2436 6739 2502 6892
rect 2628 6739 2694 6892
rect 2820 6739 2886 6892
rect 3012 6739 3078 6892
rect 3204 6739 3270 6892
rect 3688 6739 3754 6892
rect 3880 6739 3946 6892
rect 4072 6739 4138 6892
rect 4264 6739 4330 6892
rect 4456 6739 4522 6892
rect 4648 6739 4714 6892
rect 4840 6739 4906 6892
rect 5032 6739 5098 6892
rect 5516 6739 5582 6892
rect 5708 6739 5774 6892
rect 5900 6739 5966 6892
rect 6092 6739 6158 6892
rect 6284 6739 6350 6892
rect 6476 6739 6542 6892
rect 6668 6739 6734 6892
rect 6860 6739 6926 6892
rect 7344 6739 7410 6892
rect 7536 6739 7602 6892
rect 7728 6739 7794 6892
rect 7920 6739 7986 6892
rect 8112 6739 8178 6892
rect 8304 6739 8370 6892
rect 8496 6739 8562 6892
rect 8688 6739 8754 6892
rect 9172 6739 9238 6892
rect 9364 6739 9430 6892
rect 9556 6739 9622 6892
rect 9748 6739 9814 6892
rect 9940 6739 10006 6892
rect 10132 6739 10198 6892
rect 10324 6739 10390 6892
rect 10516 6739 10582 6892
rect 11000 6739 11066 6892
rect 11192 6739 11258 6892
rect 11384 6739 11450 6892
rect 11576 6739 11642 6892
rect 11768 6739 11834 6892
rect 11960 6739 12026 6892
rect 12152 6739 12218 6892
rect 12344 6739 12410 6892
rect 12828 6739 12894 6892
rect 13020 6739 13086 6892
rect 13212 6739 13278 6892
rect 13404 6739 13470 6892
rect 13596 6739 13662 6892
rect 13788 6739 13854 6892
rect 13980 6739 14046 6892
rect 14172 6739 14238 6892
rect 14656 6739 14722 6892
rect 14848 6739 14914 6892
rect 15040 6739 15106 6892
rect 15232 6739 15298 6892
rect 15424 6739 15490 6892
rect 15616 6739 15682 6892
rect 15808 6739 15874 6892
rect 16000 6739 16066 6892
rect 16484 6739 16550 6892
rect 16676 6739 16742 6892
rect 16868 6739 16934 6892
rect 17060 6739 17126 6892
rect 17252 6739 17318 6892
rect 17444 6739 17510 6892
rect 17636 6739 17702 6892
rect 17828 6739 17894 6892
rect 18312 6739 18378 6892
rect 18504 6739 18570 6892
rect 18696 6739 18762 6892
rect 18888 6739 18954 6892
rect 19080 6739 19146 6892
rect 19272 6739 19338 6892
rect 19464 6739 19530 6892
rect 19656 6739 19722 6892
rect 20140 6739 20206 6892
rect 20332 6739 20398 6892
rect 20524 6739 20590 6892
rect 20716 6739 20782 6892
rect 20908 6739 20974 6892
rect 21100 6739 21166 6892
rect 21292 6739 21358 6892
rect 21484 6739 21550 6892
rect 128 6526 194 6679
rect 320 6526 386 6679
rect 512 6526 578 6679
rect 704 6526 770 6679
rect 896 6526 962 6679
rect 1088 6526 1154 6679
rect 1280 6526 1346 6679
rect 1472 6526 1528 6679
rect 1956 6526 2022 6679
rect 2148 6526 2214 6679
rect 2340 6526 2406 6679
rect 2532 6526 2598 6679
rect 2724 6526 2790 6679
rect 2916 6526 2982 6679
rect 3108 6526 3174 6679
rect 3300 6526 3356 6679
rect 3784 6526 3850 6679
rect 3976 6526 4042 6679
rect 4168 6526 4234 6679
rect 4360 6526 4426 6679
rect 4552 6526 4618 6679
rect 4744 6526 4810 6679
rect 4936 6526 5002 6679
rect 5128 6526 5184 6679
rect 5612 6526 5678 6679
rect 5804 6526 5870 6679
rect 5996 6526 6062 6679
rect 6188 6526 6254 6679
rect 6380 6526 6446 6679
rect 6572 6526 6638 6679
rect 6764 6526 6830 6679
rect 6956 6526 7012 6679
rect 7440 6526 7506 6679
rect 7632 6526 7698 6679
rect 7824 6526 7890 6679
rect 8016 6526 8082 6679
rect 8208 6526 8274 6679
rect 8400 6526 8466 6679
rect 8592 6526 8658 6679
rect 8784 6526 8840 6679
rect 9268 6526 9334 6679
rect 9460 6526 9526 6679
rect 9652 6526 9718 6679
rect 9844 6526 9910 6679
rect 10036 6526 10102 6679
rect 10228 6526 10294 6679
rect 10420 6526 10486 6679
rect 10612 6526 10668 6679
rect 11096 6526 11162 6679
rect 11288 6526 11354 6679
rect 11480 6526 11546 6679
rect 11672 6526 11738 6679
rect 11864 6526 11930 6679
rect 12056 6526 12122 6679
rect 12248 6526 12314 6679
rect 12440 6526 12496 6679
rect 12924 6526 12990 6679
rect 13116 6526 13182 6679
rect 13308 6526 13374 6679
rect 13500 6526 13566 6679
rect 13692 6526 13758 6679
rect 13884 6526 13950 6679
rect 14076 6526 14142 6679
rect 14268 6526 14324 6679
rect 14752 6526 14818 6679
rect 14944 6526 15010 6679
rect 15136 6526 15202 6679
rect 15328 6526 15394 6679
rect 15520 6526 15586 6679
rect 15712 6526 15778 6679
rect 15904 6526 15970 6679
rect 16096 6526 16152 6679
rect 16580 6526 16646 6679
rect 16772 6526 16838 6679
rect 16964 6526 17030 6679
rect 17156 6526 17222 6679
rect 17348 6526 17414 6679
rect 17540 6526 17606 6679
rect 17732 6526 17798 6679
rect 17924 6526 17980 6679
rect 18408 6526 18474 6679
rect 18600 6526 18666 6679
rect 18792 6526 18858 6679
rect 18984 6526 19050 6679
rect 19176 6526 19242 6679
rect 19368 6526 19434 6679
rect 19560 6526 19626 6679
rect 19752 6526 19808 6679
rect 20236 6526 20302 6679
rect 20428 6526 20494 6679
rect 20620 6526 20686 6679
rect 20812 6526 20878 6679
rect 21004 6526 21070 6679
rect 21196 6526 21262 6679
rect 21388 6526 21454 6679
rect 21580 6526 21636 6679
rect 32 6025 98 6178
rect 224 6025 290 6178
rect 416 6025 482 6178
rect 608 6025 674 6178
rect 800 6025 866 6178
rect 992 6025 1058 6178
rect 1184 6025 1250 6178
rect 1376 6025 1442 6178
rect 1860 6025 1926 6178
rect 2052 6025 2118 6178
rect 2244 6025 2310 6178
rect 2436 6025 2502 6178
rect 2628 6025 2694 6178
rect 2820 6025 2886 6178
rect 3012 6025 3078 6178
rect 3204 6025 3270 6178
rect 3688 6025 3754 6178
rect 3880 6025 3946 6178
rect 4072 6025 4138 6178
rect 4264 6025 4330 6178
rect 4456 6025 4522 6178
rect 4648 6025 4714 6178
rect 4840 6025 4906 6178
rect 5032 6025 5098 6178
rect 5516 6025 5582 6178
rect 5708 6025 5774 6178
rect 5900 6025 5966 6178
rect 6092 6025 6158 6178
rect 6284 6025 6350 6178
rect 6476 6025 6542 6178
rect 6668 6025 6734 6178
rect 6860 6025 6926 6178
rect 7344 6025 7410 6178
rect 7536 6025 7602 6178
rect 7728 6025 7794 6178
rect 7920 6025 7986 6178
rect 8112 6025 8178 6178
rect 8304 6025 8370 6178
rect 8496 6025 8562 6178
rect 8688 6025 8754 6178
rect 9172 6025 9238 6178
rect 9364 6025 9430 6178
rect 9556 6025 9622 6178
rect 9748 6025 9814 6178
rect 9940 6025 10006 6178
rect 10132 6025 10198 6178
rect 10324 6025 10390 6178
rect 10516 6025 10582 6178
rect 11000 6025 11066 6178
rect 11192 6025 11258 6178
rect 11384 6025 11450 6178
rect 11576 6025 11642 6178
rect 11768 6025 11834 6178
rect 11960 6025 12026 6178
rect 12152 6025 12218 6178
rect 12344 6025 12410 6178
rect 12828 6025 12894 6178
rect 13020 6025 13086 6178
rect 13212 6025 13278 6178
rect 13404 6025 13470 6178
rect 13596 6025 13662 6178
rect 13788 6025 13854 6178
rect 13980 6025 14046 6178
rect 14172 6025 14238 6178
rect 14656 6025 14722 6178
rect 14848 6025 14914 6178
rect 15040 6025 15106 6178
rect 15232 6025 15298 6178
rect 15424 6025 15490 6178
rect 15616 6025 15682 6178
rect 15808 6025 15874 6178
rect 16000 6025 16066 6178
rect 16484 6025 16550 6178
rect 16676 6025 16742 6178
rect 16868 6025 16934 6178
rect 17060 6025 17126 6178
rect 17252 6025 17318 6178
rect 17444 6025 17510 6178
rect 17636 6025 17702 6178
rect 17828 6025 17894 6178
rect 18312 6025 18378 6178
rect 18504 6025 18570 6178
rect 18696 6025 18762 6178
rect 18888 6025 18954 6178
rect 19080 6025 19146 6178
rect 19272 6025 19338 6178
rect 19464 6025 19530 6178
rect 19656 6025 19722 6178
rect 20140 6025 20206 6178
rect 20332 6025 20398 6178
rect 20524 6025 20590 6178
rect 20716 6025 20782 6178
rect 20908 6025 20974 6178
rect 21100 6025 21166 6178
rect 21292 6025 21358 6178
rect 21484 6025 21550 6178
rect 128 5812 194 5965
rect 320 5812 386 5965
rect 512 5812 578 5965
rect 704 5812 770 5965
rect 896 5812 962 5965
rect 1088 5812 1154 5965
rect 1280 5812 1346 5965
rect 1472 5812 1528 5965
rect 1956 5812 2022 5965
rect 2148 5812 2214 5965
rect 2340 5812 2406 5965
rect 2532 5812 2598 5965
rect 2724 5812 2790 5965
rect 2916 5812 2982 5965
rect 3108 5812 3174 5965
rect 3300 5812 3356 5965
rect 3784 5812 3850 5965
rect 3976 5812 4042 5965
rect 4168 5812 4234 5965
rect 4360 5812 4426 5965
rect 4552 5812 4618 5965
rect 4744 5812 4810 5965
rect 4936 5812 5002 5965
rect 5128 5812 5184 5965
rect 5612 5812 5678 5965
rect 5804 5812 5870 5965
rect 5996 5812 6062 5965
rect 6188 5812 6254 5965
rect 6380 5812 6446 5965
rect 6572 5812 6638 5965
rect 6764 5812 6830 5965
rect 6956 5812 7012 5965
rect 7440 5812 7506 5965
rect 7632 5812 7698 5965
rect 7824 5812 7890 5965
rect 8016 5812 8082 5965
rect 8208 5812 8274 5965
rect 8400 5812 8466 5965
rect 8592 5812 8658 5965
rect 8784 5812 8840 5965
rect 9268 5812 9334 5965
rect 9460 5812 9526 5965
rect 9652 5812 9718 5965
rect 9844 5812 9910 5965
rect 10036 5812 10102 5965
rect 10228 5812 10294 5965
rect 10420 5812 10486 5965
rect 10612 5812 10668 5965
rect 11096 5812 11162 5965
rect 11288 5812 11354 5965
rect 11480 5812 11546 5965
rect 11672 5812 11738 5965
rect 11864 5812 11930 5965
rect 12056 5812 12122 5965
rect 12248 5812 12314 5965
rect 12440 5812 12496 5965
rect 12924 5812 12990 5965
rect 13116 5812 13182 5965
rect 13308 5812 13374 5965
rect 13500 5812 13566 5965
rect 13692 5812 13758 5965
rect 13884 5812 13950 5965
rect 14076 5812 14142 5965
rect 14268 5812 14324 5965
rect 14752 5812 14818 5965
rect 14944 5812 15010 5965
rect 15136 5812 15202 5965
rect 15328 5812 15394 5965
rect 15520 5812 15586 5965
rect 15712 5812 15778 5965
rect 15904 5812 15970 5965
rect 16096 5812 16152 5965
rect 16580 5812 16646 5965
rect 16772 5812 16838 5965
rect 16964 5812 17030 5965
rect 17156 5812 17222 5965
rect 17348 5812 17414 5965
rect 17540 5812 17606 5965
rect 17732 5812 17798 5965
rect 17924 5812 17980 5965
rect 18408 5812 18474 5965
rect 18600 5812 18666 5965
rect 18792 5812 18858 5965
rect 18984 5812 19050 5965
rect 19176 5812 19242 5965
rect 19368 5812 19434 5965
rect 19560 5812 19626 5965
rect 19752 5812 19808 5965
rect 20236 5812 20302 5965
rect 20428 5812 20494 5965
rect 20620 5812 20686 5965
rect 20812 5812 20878 5965
rect 21004 5812 21070 5965
rect 21196 5812 21262 5965
rect 21388 5812 21454 5965
rect 21580 5812 21636 5965
rect 32 5311 98 5464
rect 224 5311 290 5464
rect 416 5311 482 5464
rect 608 5311 674 5464
rect 800 5311 866 5464
rect 992 5311 1058 5464
rect 1184 5311 1250 5464
rect 1376 5311 1442 5464
rect 1860 5311 1926 5464
rect 2052 5311 2118 5464
rect 2244 5311 2310 5464
rect 2436 5311 2502 5464
rect 2628 5311 2694 5464
rect 2820 5311 2886 5464
rect 3012 5311 3078 5464
rect 3204 5311 3270 5464
rect 3688 5311 3754 5464
rect 3880 5311 3946 5464
rect 4072 5311 4138 5464
rect 4264 5311 4330 5464
rect 4456 5311 4522 5464
rect 4648 5311 4714 5464
rect 4840 5311 4906 5464
rect 5032 5311 5098 5464
rect 5516 5311 5582 5464
rect 5708 5311 5774 5464
rect 5900 5311 5966 5464
rect 6092 5311 6158 5464
rect 6284 5311 6350 5464
rect 6476 5311 6542 5464
rect 6668 5311 6734 5464
rect 6860 5311 6926 5464
rect 7344 5311 7410 5464
rect 7536 5311 7602 5464
rect 7728 5311 7794 5464
rect 7920 5311 7986 5464
rect 8112 5311 8178 5464
rect 8304 5311 8370 5464
rect 8496 5311 8562 5464
rect 8688 5311 8754 5464
rect 9172 5311 9238 5464
rect 9364 5311 9430 5464
rect 9556 5311 9622 5464
rect 9748 5311 9814 5464
rect 9940 5311 10006 5464
rect 10132 5311 10198 5464
rect 10324 5311 10390 5464
rect 10516 5311 10582 5464
rect 11000 5311 11066 5464
rect 11192 5311 11258 5464
rect 11384 5311 11450 5464
rect 11576 5311 11642 5464
rect 11768 5311 11834 5464
rect 11960 5311 12026 5464
rect 12152 5311 12218 5464
rect 12344 5311 12410 5464
rect 12828 5311 12894 5464
rect 13020 5311 13086 5464
rect 13212 5311 13278 5464
rect 13404 5311 13470 5464
rect 13596 5311 13662 5464
rect 13788 5311 13854 5464
rect 13980 5311 14046 5464
rect 14172 5311 14238 5464
rect 14656 5311 14722 5464
rect 14848 5311 14914 5464
rect 15040 5311 15106 5464
rect 15232 5311 15298 5464
rect 15424 5311 15490 5464
rect 15616 5311 15682 5464
rect 15808 5311 15874 5464
rect 16000 5311 16066 5464
rect 16484 5311 16550 5464
rect 16676 5311 16742 5464
rect 16868 5311 16934 5464
rect 17060 5311 17126 5464
rect 17252 5311 17318 5464
rect 17444 5311 17510 5464
rect 17636 5311 17702 5464
rect 17828 5311 17894 5464
rect 18312 5311 18378 5464
rect 18504 5311 18570 5464
rect 18696 5311 18762 5464
rect 18888 5311 18954 5464
rect 19080 5311 19146 5464
rect 19272 5311 19338 5464
rect 19464 5311 19530 5464
rect 19656 5311 19722 5464
rect 20140 5311 20206 5464
rect 20332 5311 20398 5464
rect 20524 5311 20590 5464
rect 20716 5311 20782 5464
rect 20908 5311 20974 5464
rect 21100 5311 21166 5464
rect 21292 5311 21358 5464
rect 21484 5311 21550 5464
rect 128 5098 194 5251
rect 320 5098 386 5251
rect 512 5098 578 5251
rect 704 5098 770 5251
rect 896 5098 962 5251
rect 1088 5098 1154 5251
rect 1280 5098 1346 5251
rect 1472 5098 1528 5251
rect 1956 5098 2022 5251
rect 2148 5098 2214 5251
rect 2340 5098 2406 5251
rect 2532 5098 2598 5251
rect 2724 5098 2790 5251
rect 2916 5098 2982 5251
rect 3108 5098 3174 5251
rect 3300 5098 3356 5251
rect 3784 5098 3850 5251
rect 3976 5098 4042 5251
rect 4168 5098 4234 5251
rect 4360 5098 4426 5251
rect 4552 5098 4618 5251
rect 4744 5098 4810 5251
rect 4936 5098 5002 5251
rect 5128 5098 5184 5251
rect 5612 5098 5678 5251
rect 5804 5098 5870 5251
rect 5996 5098 6062 5251
rect 6188 5098 6254 5251
rect 6380 5098 6446 5251
rect 6572 5098 6638 5251
rect 6764 5098 6830 5251
rect 6956 5098 7012 5251
rect 7440 5098 7506 5251
rect 7632 5098 7698 5251
rect 7824 5098 7890 5251
rect 8016 5098 8082 5251
rect 8208 5098 8274 5251
rect 8400 5098 8466 5251
rect 8592 5098 8658 5251
rect 8784 5098 8840 5251
rect 9268 5098 9334 5251
rect 9460 5098 9526 5251
rect 9652 5098 9718 5251
rect 9844 5098 9910 5251
rect 10036 5098 10102 5251
rect 10228 5098 10294 5251
rect 10420 5098 10486 5251
rect 10612 5098 10668 5251
rect 11096 5098 11162 5251
rect 11288 5098 11354 5251
rect 11480 5098 11546 5251
rect 11672 5098 11738 5251
rect 11864 5098 11930 5251
rect 12056 5098 12122 5251
rect 12248 5098 12314 5251
rect 12440 5098 12496 5251
rect 12924 5098 12990 5251
rect 13116 5098 13182 5251
rect 13308 5098 13374 5251
rect 13500 5098 13566 5251
rect 13692 5098 13758 5251
rect 13884 5098 13950 5251
rect 14076 5098 14142 5251
rect 14268 5098 14324 5251
rect 14752 5098 14818 5251
rect 14944 5098 15010 5251
rect 15136 5098 15202 5251
rect 15328 5098 15394 5251
rect 15520 5098 15586 5251
rect 15712 5098 15778 5251
rect 15904 5098 15970 5251
rect 16096 5098 16152 5251
rect 16580 5098 16646 5251
rect 16772 5098 16838 5251
rect 16964 5098 17030 5251
rect 17156 5098 17222 5251
rect 17348 5098 17414 5251
rect 17540 5098 17606 5251
rect 17732 5098 17798 5251
rect 17924 5098 17980 5251
rect 18408 5098 18474 5251
rect 18600 5098 18666 5251
rect 18792 5098 18858 5251
rect 18984 5098 19050 5251
rect 19176 5098 19242 5251
rect 19368 5098 19434 5251
rect 19560 5098 19626 5251
rect 19752 5098 19808 5251
rect 20236 5098 20302 5251
rect 20428 5098 20494 5251
rect 20620 5098 20686 5251
rect 20812 5098 20878 5251
rect 21004 5098 21070 5251
rect 21196 5098 21262 5251
rect 21388 5098 21454 5251
rect 21580 5098 21636 5251
rect 32 4597 98 4750
rect 224 4597 290 4750
rect 416 4597 482 4750
rect 608 4597 674 4750
rect 800 4597 866 4750
rect 992 4597 1058 4750
rect 1184 4597 1250 4750
rect 1376 4597 1442 4750
rect 1860 4597 1926 4750
rect 2052 4597 2118 4750
rect 2244 4597 2310 4750
rect 2436 4597 2502 4750
rect 2628 4597 2694 4750
rect 2820 4597 2886 4750
rect 3012 4597 3078 4750
rect 3204 4597 3270 4750
rect 3688 4597 3754 4750
rect 3880 4597 3946 4750
rect 4072 4597 4138 4750
rect 4264 4597 4330 4750
rect 4456 4597 4522 4750
rect 4648 4597 4714 4750
rect 4840 4597 4906 4750
rect 5032 4597 5098 4750
rect 5516 4597 5582 4750
rect 5708 4597 5774 4750
rect 5900 4597 5966 4750
rect 6092 4597 6158 4750
rect 6284 4597 6350 4750
rect 6476 4597 6542 4750
rect 6668 4597 6734 4750
rect 6860 4597 6926 4750
rect 7344 4597 7410 4750
rect 7536 4597 7602 4750
rect 7728 4597 7794 4750
rect 7920 4597 7986 4750
rect 8112 4597 8178 4750
rect 8304 4597 8370 4750
rect 8496 4597 8562 4750
rect 8688 4597 8754 4750
rect 9172 4597 9238 4750
rect 9364 4597 9430 4750
rect 9556 4597 9622 4750
rect 9748 4597 9814 4750
rect 9940 4597 10006 4750
rect 10132 4597 10198 4750
rect 10324 4597 10390 4750
rect 10516 4597 10582 4750
rect 11000 4597 11066 4750
rect 11192 4597 11258 4750
rect 11384 4597 11450 4750
rect 11576 4597 11642 4750
rect 11768 4597 11834 4750
rect 11960 4597 12026 4750
rect 12152 4597 12218 4750
rect 12344 4597 12410 4750
rect 12828 4597 12894 4750
rect 13020 4597 13086 4750
rect 13212 4597 13278 4750
rect 13404 4597 13470 4750
rect 13596 4597 13662 4750
rect 13788 4597 13854 4750
rect 13980 4597 14046 4750
rect 14172 4597 14238 4750
rect 14656 4597 14722 4750
rect 14848 4597 14914 4750
rect 15040 4597 15106 4750
rect 15232 4597 15298 4750
rect 15424 4597 15490 4750
rect 15616 4597 15682 4750
rect 15808 4597 15874 4750
rect 16000 4597 16066 4750
rect 16484 4597 16550 4750
rect 16676 4597 16742 4750
rect 16868 4597 16934 4750
rect 17060 4597 17126 4750
rect 17252 4597 17318 4750
rect 17444 4597 17510 4750
rect 17636 4597 17702 4750
rect 17828 4597 17894 4750
rect 18312 4597 18378 4750
rect 18504 4597 18570 4750
rect 18696 4597 18762 4750
rect 18888 4597 18954 4750
rect 19080 4597 19146 4750
rect 19272 4597 19338 4750
rect 19464 4597 19530 4750
rect 19656 4597 19722 4750
rect 20140 4597 20206 4750
rect 20332 4597 20398 4750
rect 20524 4597 20590 4750
rect 20716 4597 20782 4750
rect 20908 4597 20974 4750
rect 21100 4597 21166 4750
rect 21292 4597 21358 4750
rect 21484 4597 21550 4750
rect 128 4384 194 4537
rect 320 4384 386 4537
rect 512 4384 578 4537
rect 704 4384 770 4537
rect 896 4384 962 4537
rect 1088 4384 1154 4537
rect 1280 4384 1346 4537
rect 1472 4384 1528 4537
rect 1956 4384 2022 4537
rect 2148 4384 2214 4537
rect 2340 4384 2406 4537
rect 2532 4384 2598 4537
rect 2724 4384 2790 4537
rect 2916 4384 2982 4537
rect 3108 4384 3174 4537
rect 3300 4384 3356 4537
rect 3784 4384 3850 4537
rect 3976 4384 4042 4537
rect 4168 4384 4234 4537
rect 4360 4384 4426 4537
rect 4552 4384 4618 4537
rect 4744 4384 4810 4537
rect 4936 4384 5002 4537
rect 5128 4384 5184 4537
rect 5612 4384 5678 4537
rect 5804 4384 5870 4537
rect 5996 4384 6062 4537
rect 6188 4384 6254 4537
rect 6380 4384 6446 4537
rect 6572 4384 6638 4537
rect 6764 4384 6830 4537
rect 6956 4384 7012 4537
rect 7440 4384 7506 4537
rect 7632 4384 7698 4537
rect 7824 4384 7890 4537
rect 8016 4384 8082 4537
rect 8208 4384 8274 4537
rect 8400 4384 8466 4537
rect 8592 4384 8658 4537
rect 8784 4384 8840 4537
rect 9268 4384 9334 4537
rect 9460 4384 9526 4537
rect 9652 4384 9718 4537
rect 9844 4384 9910 4537
rect 10036 4384 10102 4537
rect 10228 4384 10294 4537
rect 10420 4384 10486 4537
rect 10612 4384 10668 4537
rect 11096 4384 11162 4537
rect 11288 4384 11354 4537
rect 11480 4384 11546 4537
rect 11672 4384 11738 4537
rect 11864 4384 11930 4537
rect 12056 4384 12122 4537
rect 12248 4384 12314 4537
rect 12440 4384 12496 4537
rect 12924 4384 12990 4537
rect 13116 4384 13182 4537
rect 13308 4384 13374 4537
rect 13500 4384 13566 4537
rect 13692 4384 13758 4537
rect 13884 4384 13950 4537
rect 14076 4384 14142 4537
rect 14268 4384 14324 4537
rect 14752 4384 14818 4537
rect 14944 4384 15010 4537
rect 15136 4384 15202 4537
rect 15328 4384 15394 4537
rect 15520 4384 15586 4537
rect 15712 4384 15778 4537
rect 15904 4384 15970 4537
rect 16096 4384 16152 4537
rect 16580 4384 16646 4537
rect 16772 4384 16838 4537
rect 16964 4384 17030 4537
rect 17156 4384 17222 4537
rect 17348 4384 17414 4537
rect 17540 4384 17606 4537
rect 17732 4384 17798 4537
rect 17924 4384 17980 4537
rect 18408 4384 18474 4537
rect 18600 4384 18666 4537
rect 18792 4384 18858 4537
rect 18984 4384 19050 4537
rect 19176 4384 19242 4537
rect 19368 4384 19434 4537
rect 19560 4384 19626 4537
rect 19752 4384 19808 4537
rect 20236 4384 20302 4537
rect 20428 4384 20494 4537
rect 20620 4384 20686 4537
rect 20812 4384 20878 4537
rect 21004 4384 21070 4537
rect 21196 4384 21262 4537
rect 21388 4384 21454 4537
rect 21580 4384 21636 4537
rect 32 3883 98 4036
rect 224 3883 290 4036
rect 416 3883 482 4036
rect 608 3883 674 4036
rect 800 3883 866 4036
rect 992 3883 1058 4036
rect 1184 3883 1250 4036
rect 1376 3883 1442 4036
rect 1860 3883 1926 4036
rect 2052 3883 2118 4036
rect 2244 3883 2310 4036
rect 2436 3883 2502 4036
rect 2628 3883 2694 4036
rect 2820 3883 2886 4036
rect 3012 3883 3078 4036
rect 3204 3883 3270 4036
rect 3688 3883 3754 4036
rect 3880 3883 3946 4036
rect 4072 3883 4138 4036
rect 4264 3883 4330 4036
rect 4456 3883 4522 4036
rect 4648 3883 4714 4036
rect 4840 3883 4906 4036
rect 5032 3883 5098 4036
rect 5516 3883 5582 4036
rect 5708 3883 5774 4036
rect 5900 3883 5966 4036
rect 6092 3883 6158 4036
rect 6284 3883 6350 4036
rect 6476 3883 6542 4036
rect 6668 3883 6734 4036
rect 6860 3883 6926 4036
rect 7344 3883 7410 4036
rect 7536 3883 7602 4036
rect 7728 3883 7794 4036
rect 7920 3883 7986 4036
rect 8112 3883 8178 4036
rect 8304 3883 8370 4036
rect 8496 3883 8562 4036
rect 8688 3883 8754 4036
rect 9172 3883 9238 4036
rect 9364 3883 9430 4036
rect 9556 3883 9622 4036
rect 9748 3883 9814 4036
rect 9940 3883 10006 4036
rect 10132 3883 10198 4036
rect 10324 3883 10390 4036
rect 10516 3883 10582 4036
rect 11000 3883 11066 4036
rect 11192 3883 11258 4036
rect 11384 3883 11450 4036
rect 11576 3883 11642 4036
rect 11768 3883 11834 4036
rect 11960 3883 12026 4036
rect 12152 3883 12218 4036
rect 12344 3883 12410 4036
rect 12828 3883 12894 4036
rect 13020 3883 13086 4036
rect 13212 3883 13278 4036
rect 13404 3883 13470 4036
rect 13596 3883 13662 4036
rect 13788 3883 13854 4036
rect 13980 3883 14046 4036
rect 14172 3883 14238 4036
rect 14656 3883 14722 4036
rect 14848 3883 14914 4036
rect 15040 3883 15106 4036
rect 15232 3883 15298 4036
rect 15424 3883 15490 4036
rect 15616 3883 15682 4036
rect 15808 3883 15874 4036
rect 16000 3883 16066 4036
rect 16484 3883 16550 4036
rect 16676 3883 16742 4036
rect 16868 3883 16934 4036
rect 17060 3883 17126 4036
rect 17252 3883 17318 4036
rect 17444 3883 17510 4036
rect 17636 3883 17702 4036
rect 17828 3883 17894 4036
rect 18312 3883 18378 4036
rect 18504 3883 18570 4036
rect 18696 3883 18762 4036
rect 18888 3883 18954 4036
rect 19080 3883 19146 4036
rect 19272 3883 19338 4036
rect 19464 3883 19530 4036
rect 19656 3883 19722 4036
rect 20140 3883 20206 4036
rect 20332 3883 20398 4036
rect 20524 3883 20590 4036
rect 20716 3883 20782 4036
rect 20908 3883 20974 4036
rect 21100 3883 21166 4036
rect 21292 3883 21358 4036
rect 21484 3883 21550 4036
rect 128 3670 194 3823
rect 320 3670 386 3823
rect 512 3670 578 3823
rect 704 3670 770 3823
rect 896 3670 962 3823
rect 1088 3670 1154 3823
rect 1280 3670 1346 3823
rect 1472 3670 1528 3823
rect 1956 3670 2022 3823
rect 2148 3670 2214 3823
rect 2340 3670 2406 3823
rect 2532 3670 2598 3823
rect 2724 3670 2790 3823
rect 2916 3670 2982 3823
rect 3108 3670 3174 3823
rect 3300 3670 3356 3823
rect 3784 3670 3850 3823
rect 3976 3670 4042 3823
rect 4168 3670 4234 3823
rect 4360 3670 4426 3823
rect 4552 3670 4618 3823
rect 4744 3670 4810 3823
rect 4936 3670 5002 3823
rect 5128 3670 5184 3823
rect 5612 3670 5678 3823
rect 5804 3670 5870 3823
rect 5996 3670 6062 3823
rect 6188 3670 6254 3823
rect 6380 3670 6446 3823
rect 6572 3670 6638 3823
rect 6764 3670 6830 3823
rect 6956 3670 7012 3823
rect 7440 3670 7506 3823
rect 7632 3670 7698 3823
rect 7824 3670 7890 3823
rect 8016 3670 8082 3823
rect 8208 3670 8274 3823
rect 8400 3670 8466 3823
rect 8592 3670 8658 3823
rect 8784 3670 8840 3823
rect 9268 3670 9334 3823
rect 9460 3670 9526 3823
rect 9652 3670 9718 3823
rect 9844 3670 9910 3823
rect 10036 3670 10102 3823
rect 10228 3670 10294 3823
rect 10420 3670 10486 3823
rect 10612 3670 10668 3823
rect 11096 3670 11162 3823
rect 11288 3670 11354 3823
rect 11480 3670 11546 3823
rect 11672 3670 11738 3823
rect 11864 3670 11930 3823
rect 12056 3670 12122 3823
rect 12248 3670 12314 3823
rect 12440 3670 12496 3823
rect 12924 3670 12990 3823
rect 13116 3670 13182 3823
rect 13308 3670 13374 3823
rect 13500 3670 13566 3823
rect 13692 3670 13758 3823
rect 13884 3670 13950 3823
rect 14076 3670 14142 3823
rect 14268 3670 14324 3823
rect 14752 3670 14818 3823
rect 14944 3670 15010 3823
rect 15136 3670 15202 3823
rect 15328 3670 15394 3823
rect 15520 3670 15586 3823
rect 15712 3670 15778 3823
rect 15904 3670 15970 3823
rect 16096 3670 16152 3823
rect 16580 3670 16646 3823
rect 16772 3670 16838 3823
rect 16964 3670 17030 3823
rect 17156 3670 17222 3823
rect 17348 3670 17414 3823
rect 17540 3670 17606 3823
rect 17732 3670 17798 3823
rect 17924 3670 17980 3823
rect 18408 3670 18474 3823
rect 18600 3670 18666 3823
rect 18792 3670 18858 3823
rect 18984 3670 19050 3823
rect 19176 3670 19242 3823
rect 19368 3670 19434 3823
rect 19560 3670 19626 3823
rect 19752 3670 19808 3823
rect 20236 3670 20302 3823
rect 20428 3670 20494 3823
rect 20620 3670 20686 3823
rect 20812 3670 20878 3823
rect 21004 3670 21070 3823
rect 21196 3670 21262 3823
rect 21388 3670 21454 3823
rect 21580 3670 21636 3823
rect 32 3169 98 3322
rect 224 3169 290 3322
rect 416 3169 482 3322
rect 608 3169 674 3322
rect 800 3169 866 3322
rect 992 3169 1058 3322
rect 1184 3169 1250 3322
rect 1376 3169 1442 3322
rect 1860 3169 1926 3322
rect 2052 3169 2118 3322
rect 2244 3169 2310 3322
rect 2436 3169 2502 3322
rect 2628 3169 2694 3322
rect 2820 3169 2886 3322
rect 3012 3169 3078 3322
rect 3204 3169 3270 3322
rect 3688 3169 3754 3322
rect 3880 3169 3946 3322
rect 4072 3169 4138 3322
rect 4264 3169 4330 3322
rect 4456 3169 4522 3322
rect 4648 3169 4714 3322
rect 4840 3169 4906 3322
rect 5032 3169 5098 3322
rect 5516 3169 5582 3322
rect 5708 3169 5774 3322
rect 5900 3169 5966 3322
rect 6092 3169 6158 3322
rect 6284 3169 6350 3322
rect 6476 3169 6542 3322
rect 6668 3169 6734 3322
rect 6860 3169 6926 3322
rect 7344 3169 7410 3322
rect 7536 3169 7602 3322
rect 7728 3169 7794 3322
rect 7920 3169 7986 3322
rect 8112 3169 8178 3322
rect 8304 3169 8370 3322
rect 8496 3169 8562 3322
rect 8688 3169 8754 3322
rect 9172 3169 9238 3322
rect 9364 3169 9430 3322
rect 9556 3169 9622 3322
rect 9748 3169 9814 3322
rect 9940 3169 10006 3322
rect 10132 3169 10198 3322
rect 10324 3169 10390 3322
rect 10516 3169 10582 3322
rect 11000 3169 11066 3322
rect 11192 3169 11258 3322
rect 11384 3169 11450 3322
rect 11576 3169 11642 3322
rect 11768 3169 11834 3322
rect 11960 3169 12026 3322
rect 12152 3169 12218 3322
rect 12344 3169 12410 3322
rect 12828 3169 12894 3322
rect 13020 3169 13086 3322
rect 13212 3169 13278 3322
rect 13404 3169 13470 3322
rect 13596 3169 13662 3322
rect 13788 3169 13854 3322
rect 13980 3169 14046 3322
rect 14172 3169 14238 3322
rect 14656 3169 14722 3322
rect 14848 3169 14914 3322
rect 15040 3169 15106 3322
rect 15232 3169 15298 3322
rect 15424 3169 15490 3322
rect 15616 3169 15682 3322
rect 15808 3169 15874 3322
rect 16000 3169 16066 3322
rect 16484 3169 16550 3322
rect 16676 3169 16742 3322
rect 16868 3169 16934 3322
rect 17060 3169 17126 3322
rect 17252 3169 17318 3322
rect 17444 3169 17510 3322
rect 17636 3169 17702 3322
rect 17828 3169 17894 3322
rect 18312 3169 18378 3322
rect 18504 3169 18570 3322
rect 18696 3169 18762 3322
rect 18888 3169 18954 3322
rect 19080 3169 19146 3322
rect 19272 3169 19338 3322
rect 19464 3169 19530 3322
rect 19656 3169 19722 3322
rect 20140 3169 20206 3322
rect 20332 3169 20398 3322
rect 20524 3169 20590 3322
rect 20716 3169 20782 3322
rect 20908 3169 20974 3322
rect 21100 3169 21166 3322
rect 21292 3169 21358 3322
rect 21484 3169 21550 3322
rect 128 2956 194 3109
rect 320 2956 386 3109
rect 512 2956 578 3109
rect 704 2956 770 3109
rect 896 2956 962 3109
rect 1088 2956 1154 3109
rect 1280 2956 1346 3109
rect 1472 2956 1528 3109
rect 1956 2956 2022 3109
rect 2148 2956 2214 3109
rect 2340 2956 2406 3109
rect 2532 2956 2598 3109
rect 2724 2956 2790 3109
rect 2916 2956 2982 3109
rect 3108 2956 3174 3109
rect 3300 2956 3356 3109
rect 3784 2956 3850 3109
rect 3976 2956 4042 3109
rect 4168 2956 4234 3109
rect 4360 2956 4426 3109
rect 4552 2956 4618 3109
rect 4744 2956 4810 3109
rect 4936 2956 5002 3109
rect 5128 2956 5184 3109
rect 5612 2956 5678 3109
rect 5804 2956 5870 3109
rect 5996 2956 6062 3109
rect 6188 2956 6254 3109
rect 6380 2956 6446 3109
rect 6572 2956 6638 3109
rect 6764 2956 6830 3109
rect 6956 2956 7012 3109
rect 7440 2956 7506 3109
rect 7632 2956 7698 3109
rect 7824 2956 7890 3109
rect 8016 2956 8082 3109
rect 8208 2956 8274 3109
rect 8400 2956 8466 3109
rect 8592 2956 8658 3109
rect 8784 2956 8840 3109
rect 9268 2956 9334 3109
rect 9460 2956 9526 3109
rect 9652 2956 9718 3109
rect 9844 2956 9910 3109
rect 10036 2956 10102 3109
rect 10228 2956 10294 3109
rect 10420 2956 10486 3109
rect 10612 2956 10668 3109
rect 11096 2956 11162 3109
rect 11288 2956 11354 3109
rect 11480 2956 11546 3109
rect 11672 2956 11738 3109
rect 11864 2956 11930 3109
rect 12056 2956 12122 3109
rect 12248 2956 12314 3109
rect 12440 2956 12496 3109
rect 12924 2956 12990 3109
rect 13116 2956 13182 3109
rect 13308 2956 13374 3109
rect 13500 2956 13566 3109
rect 13692 2956 13758 3109
rect 13884 2956 13950 3109
rect 14076 2956 14142 3109
rect 14268 2956 14324 3109
rect 14752 2956 14818 3109
rect 14944 2956 15010 3109
rect 15136 2956 15202 3109
rect 15328 2956 15394 3109
rect 15520 2956 15586 3109
rect 15712 2956 15778 3109
rect 15904 2956 15970 3109
rect 16096 2956 16152 3109
rect 16580 2956 16646 3109
rect 16772 2956 16838 3109
rect 16964 2956 17030 3109
rect 17156 2956 17222 3109
rect 17348 2956 17414 3109
rect 17540 2956 17606 3109
rect 17732 2956 17798 3109
rect 17924 2956 17980 3109
rect 18408 2956 18474 3109
rect 18600 2956 18666 3109
rect 18792 2956 18858 3109
rect 18984 2956 19050 3109
rect 19176 2956 19242 3109
rect 19368 2956 19434 3109
rect 19560 2956 19626 3109
rect 19752 2956 19808 3109
rect 20236 2956 20302 3109
rect 20428 2956 20494 3109
rect 20620 2956 20686 3109
rect 20812 2956 20878 3109
rect 21004 2956 21070 3109
rect 21196 2956 21262 3109
rect 21388 2956 21454 3109
rect 21580 2956 21636 3109
rect 32 2455 98 2608
rect 224 2455 290 2608
rect 416 2455 482 2608
rect 608 2455 674 2608
rect 800 2455 866 2608
rect 992 2455 1058 2608
rect 1184 2455 1250 2608
rect 1376 2455 1442 2608
rect 1860 2455 1926 2608
rect 2052 2455 2118 2608
rect 2244 2455 2310 2608
rect 2436 2455 2502 2608
rect 2628 2455 2694 2608
rect 2820 2455 2886 2608
rect 3012 2455 3078 2608
rect 3204 2455 3270 2608
rect 3688 2455 3754 2608
rect 3880 2455 3946 2608
rect 4072 2455 4138 2608
rect 4264 2455 4330 2608
rect 4456 2455 4522 2608
rect 4648 2455 4714 2608
rect 4840 2455 4906 2608
rect 5032 2455 5098 2608
rect 5516 2455 5582 2608
rect 5708 2455 5774 2608
rect 5900 2455 5966 2608
rect 6092 2455 6158 2608
rect 6284 2455 6350 2608
rect 6476 2455 6542 2608
rect 6668 2455 6734 2608
rect 6860 2455 6926 2608
rect 7344 2455 7410 2608
rect 7536 2455 7602 2608
rect 7728 2455 7794 2608
rect 7920 2455 7986 2608
rect 8112 2455 8178 2608
rect 8304 2455 8370 2608
rect 8496 2455 8562 2608
rect 8688 2455 8754 2608
rect 9172 2455 9238 2608
rect 9364 2455 9430 2608
rect 9556 2455 9622 2608
rect 9748 2455 9814 2608
rect 9940 2455 10006 2608
rect 10132 2455 10198 2608
rect 10324 2455 10390 2608
rect 10516 2455 10582 2608
rect 11000 2455 11066 2608
rect 11192 2455 11258 2608
rect 11384 2455 11450 2608
rect 11576 2455 11642 2608
rect 11768 2455 11834 2608
rect 11960 2455 12026 2608
rect 12152 2455 12218 2608
rect 12344 2455 12410 2608
rect 12828 2455 12894 2608
rect 13020 2455 13086 2608
rect 13212 2455 13278 2608
rect 13404 2455 13470 2608
rect 13596 2455 13662 2608
rect 13788 2455 13854 2608
rect 13980 2455 14046 2608
rect 14172 2455 14238 2608
rect 14656 2455 14722 2608
rect 14848 2455 14914 2608
rect 15040 2455 15106 2608
rect 15232 2455 15298 2608
rect 15424 2455 15490 2608
rect 15616 2455 15682 2608
rect 15808 2455 15874 2608
rect 16000 2455 16066 2608
rect 16484 2455 16550 2608
rect 16676 2455 16742 2608
rect 16868 2455 16934 2608
rect 17060 2455 17126 2608
rect 17252 2455 17318 2608
rect 17444 2455 17510 2608
rect 17636 2455 17702 2608
rect 17828 2455 17894 2608
rect 18312 2455 18378 2608
rect 18504 2455 18570 2608
rect 18696 2455 18762 2608
rect 18888 2455 18954 2608
rect 19080 2455 19146 2608
rect 19272 2455 19338 2608
rect 19464 2455 19530 2608
rect 19656 2455 19722 2608
rect 20140 2455 20206 2608
rect 20332 2455 20398 2608
rect 20524 2455 20590 2608
rect 20716 2455 20782 2608
rect 20908 2455 20974 2608
rect 21100 2455 21166 2608
rect 21292 2455 21358 2608
rect 21484 2455 21550 2608
rect 128 2242 194 2395
rect 320 2242 386 2395
rect 512 2242 578 2395
rect 704 2242 770 2395
rect 896 2242 962 2395
rect 1088 2242 1154 2395
rect 1280 2242 1346 2395
rect 1472 2242 1528 2395
rect 1956 2242 2022 2395
rect 2148 2242 2214 2395
rect 2340 2242 2406 2395
rect 2532 2242 2598 2395
rect 2724 2242 2790 2395
rect 2916 2242 2982 2395
rect 3108 2242 3174 2395
rect 3300 2242 3356 2395
rect 3784 2242 3850 2395
rect 3976 2242 4042 2395
rect 4168 2242 4234 2395
rect 4360 2242 4426 2395
rect 4552 2242 4618 2395
rect 4744 2242 4810 2395
rect 4936 2242 5002 2395
rect 5128 2242 5184 2395
rect 5612 2242 5678 2395
rect 5804 2242 5870 2395
rect 5996 2242 6062 2395
rect 6188 2242 6254 2395
rect 6380 2242 6446 2395
rect 6572 2242 6638 2395
rect 6764 2242 6830 2395
rect 6956 2242 7012 2395
rect 7440 2242 7506 2395
rect 7632 2242 7698 2395
rect 7824 2242 7890 2395
rect 8016 2242 8082 2395
rect 8208 2242 8274 2395
rect 8400 2242 8466 2395
rect 8592 2242 8658 2395
rect 8784 2242 8840 2395
rect 9268 2242 9334 2395
rect 9460 2242 9526 2395
rect 9652 2242 9718 2395
rect 9844 2242 9910 2395
rect 10036 2242 10102 2395
rect 10228 2242 10294 2395
rect 10420 2242 10486 2395
rect 10612 2242 10668 2395
rect 11096 2242 11162 2395
rect 11288 2242 11354 2395
rect 11480 2242 11546 2395
rect 11672 2242 11738 2395
rect 11864 2242 11930 2395
rect 12056 2242 12122 2395
rect 12248 2242 12314 2395
rect 12440 2242 12496 2395
rect 12924 2242 12990 2395
rect 13116 2242 13182 2395
rect 13308 2242 13374 2395
rect 13500 2242 13566 2395
rect 13692 2242 13758 2395
rect 13884 2242 13950 2395
rect 14076 2242 14142 2395
rect 14268 2242 14324 2395
rect 14752 2242 14818 2395
rect 14944 2242 15010 2395
rect 15136 2242 15202 2395
rect 15328 2242 15394 2395
rect 15520 2242 15586 2395
rect 15712 2242 15778 2395
rect 15904 2242 15970 2395
rect 16096 2242 16152 2395
rect 16580 2242 16646 2395
rect 16772 2242 16838 2395
rect 16964 2242 17030 2395
rect 17156 2242 17222 2395
rect 17348 2242 17414 2395
rect 17540 2242 17606 2395
rect 17732 2242 17798 2395
rect 17924 2242 17980 2395
rect 18408 2242 18474 2395
rect 18600 2242 18666 2395
rect 18792 2242 18858 2395
rect 18984 2242 19050 2395
rect 19176 2242 19242 2395
rect 19368 2242 19434 2395
rect 19560 2242 19626 2395
rect 19752 2242 19808 2395
rect 20236 2242 20302 2395
rect 20428 2242 20494 2395
rect 20620 2242 20686 2395
rect 20812 2242 20878 2395
rect 21004 2242 21070 2395
rect 21196 2242 21262 2395
rect 21388 2242 21454 2395
rect 21580 2242 21636 2395
rect 32 1741 98 1894
rect 224 1741 290 1894
rect 416 1741 482 1894
rect 608 1741 674 1894
rect 800 1741 866 1894
rect 992 1741 1058 1894
rect 1184 1741 1250 1894
rect 1376 1741 1442 1894
rect 1860 1741 1926 1894
rect 2052 1741 2118 1894
rect 2244 1741 2310 1894
rect 2436 1741 2502 1894
rect 2628 1741 2694 1894
rect 2820 1741 2886 1894
rect 3012 1741 3078 1894
rect 3204 1741 3270 1894
rect 3688 1741 3754 1894
rect 3880 1741 3946 1894
rect 4072 1741 4138 1894
rect 4264 1741 4330 1894
rect 4456 1741 4522 1894
rect 4648 1741 4714 1894
rect 4840 1741 4906 1894
rect 5032 1741 5098 1894
rect 5516 1741 5582 1894
rect 5708 1741 5774 1894
rect 5900 1741 5966 1894
rect 6092 1741 6158 1894
rect 6284 1741 6350 1894
rect 6476 1741 6542 1894
rect 6668 1741 6734 1894
rect 6860 1741 6926 1894
rect 7344 1741 7410 1894
rect 7536 1741 7602 1894
rect 7728 1741 7794 1894
rect 7920 1741 7986 1894
rect 8112 1741 8178 1894
rect 8304 1741 8370 1894
rect 8496 1741 8562 1894
rect 8688 1741 8754 1894
rect 9172 1741 9238 1894
rect 9364 1741 9430 1894
rect 9556 1741 9622 1894
rect 9748 1741 9814 1894
rect 9940 1741 10006 1894
rect 10132 1741 10198 1894
rect 10324 1741 10390 1894
rect 10516 1741 10582 1894
rect 11000 1741 11066 1894
rect 11192 1741 11258 1894
rect 11384 1741 11450 1894
rect 11576 1741 11642 1894
rect 11768 1741 11834 1894
rect 11960 1741 12026 1894
rect 12152 1741 12218 1894
rect 12344 1741 12410 1894
rect 12828 1741 12894 1894
rect 13020 1741 13086 1894
rect 13212 1741 13278 1894
rect 13404 1741 13470 1894
rect 13596 1741 13662 1894
rect 13788 1741 13854 1894
rect 13980 1741 14046 1894
rect 14172 1741 14238 1894
rect 14656 1741 14722 1894
rect 14848 1741 14914 1894
rect 15040 1741 15106 1894
rect 15232 1741 15298 1894
rect 15424 1741 15490 1894
rect 15616 1741 15682 1894
rect 15808 1741 15874 1894
rect 16000 1741 16066 1894
rect 16484 1741 16550 1894
rect 16676 1741 16742 1894
rect 16868 1741 16934 1894
rect 17060 1741 17126 1894
rect 17252 1741 17318 1894
rect 17444 1741 17510 1894
rect 17636 1741 17702 1894
rect 17828 1741 17894 1894
rect 18312 1741 18378 1894
rect 18504 1741 18570 1894
rect 18696 1741 18762 1894
rect 18888 1741 18954 1894
rect 19080 1741 19146 1894
rect 19272 1741 19338 1894
rect 19464 1741 19530 1894
rect 19656 1741 19722 1894
rect 20140 1741 20206 1894
rect 20332 1741 20398 1894
rect 20524 1741 20590 1894
rect 20716 1741 20782 1894
rect 20908 1741 20974 1894
rect 21100 1741 21166 1894
rect 21292 1741 21358 1894
rect 21484 1741 21550 1894
rect 128 1528 194 1681
rect 320 1528 386 1681
rect 512 1528 578 1681
rect 704 1528 770 1681
rect 896 1528 962 1681
rect 1088 1528 1154 1681
rect 1280 1528 1346 1681
rect 1472 1528 1528 1681
rect 1956 1528 2022 1681
rect 2148 1528 2214 1681
rect 2340 1528 2406 1681
rect 2532 1528 2598 1681
rect 2724 1528 2790 1681
rect 2916 1528 2982 1681
rect 3108 1528 3174 1681
rect 3300 1528 3356 1681
rect 3784 1528 3850 1681
rect 3976 1528 4042 1681
rect 4168 1528 4234 1681
rect 4360 1528 4426 1681
rect 4552 1528 4618 1681
rect 4744 1528 4810 1681
rect 4936 1528 5002 1681
rect 5128 1528 5184 1681
rect 5612 1528 5678 1681
rect 5804 1528 5870 1681
rect 5996 1528 6062 1681
rect 6188 1528 6254 1681
rect 6380 1528 6446 1681
rect 6572 1528 6638 1681
rect 6764 1528 6830 1681
rect 6956 1528 7012 1681
rect 7440 1528 7506 1681
rect 7632 1528 7698 1681
rect 7824 1528 7890 1681
rect 8016 1528 8082 1681
rect 8208 1528 8274 1681
rect 8400 1528 8466 1681
rect 8592 1528 8658 1681
rect 8784 1528 8840 1681
rect 9268 1528 9334 1681
rect 9460 1528 9526 1681
rect 9652 1528 9718 1681
rect 9844 1528 9910 1681
rect 10036 1528 10102 1681
rect 10228 1528 10294 1681
rect 10420 1528 10486 1681
rect 10612 1528 10668 1681
rect 11096 1528 11162 1681
rect 11288 1528 11354 1681
rect 11480 1528 11546 1681
rect 11672 1528 11738 1681
rect 11864 1528 11930 1681
rect 12056 1528 12122 1681
rect 12248 1528 12314 1681
rect 12440 1528 12496 1681
rect 12924 1528 12990 1681
rect 13116 1528 13182 1681
rect 13308 1528 13374 1681
rect 13500 1528 13566 1681
rect 13692 1528 13758 1681
rect 13884 1528 13950 1681
rect 14076 1528 14142 1681
rect 14268 1528 14324 1681
rect 14752 1528 14818 1681
rect 14944 1528 15010 1681
rect 15136 1528 15202 1681
rect 15328 1528 15394 1681
rect 15520 1528 15586 1681
rect 15712 1528 15778 1681
rect 15904 1528 15970 1681
rect 16096 1528 16152 1681
rect 16580 1528 16646 1681
rect 16772 1528 16838 1681
rect 16964 1528 17030 1681
rect 17156 1528 17222 1681
rect 17348 1528 17414 1681
rect 17540 1528 17606 1681
rect 17732 1528 17798 1681
rect 17924 1528 17980 1681
rect 18408 1528 18474 1681
rect 18600 1528 18666 1681
rect 18792 1528 18858 1681
rect 18984 1528 19050 1681
rect 19176 1528 19242 1681
rect 19368 1528 19434 1681
rect 19560 1528 19626 1681
rect 19752 1528 19808 1681
rect 20236 1528 20302 1681
rect 20428 1528 20494 1681
rect 20620 1528 20686 1681
rect 20812 1528 20878 1681
rect 21004 1528 21070 1681
rect 21196 1528 21262 1681
rect 21388 1528 21454 1681
rect 21580 1528 21636 1681
rect 32 1027 98 1180
rect 224 1027 290 1180
rect 416 1027 482 1180
rect 608 1027 674 1180
rect 800 1027 866 1180
rect 992 1027 1058 1180
rect 1184 1027 1250 1180
rect 1376 1027 1442 1180
rect 1860 1027 1926 1180
rect 2052 1027 2118 1180
rect 2244 1027 2310 1180
rect 2436 1027 2502 1180
rect 2628 1027 2694 1180
rect 2820 1027 2886 1180
rect 3012 1027 3078 1180
rect 3204 1027 3270 1180
rect 3688 1027 3754 1180
rect 3880 1027 3946 1180
rect 4072 1027 4138 1180
rect 4264 1027 4330 1180
rect 4456 1027 4522 1180
rect 4648 1027 4714 1180
rect 4840 1027 4906 1180
rect 5032 1027 5098 1180
rect 5516 1027 5582 1180
rect 5708 1027 5774 1180
rect 5900 1027 5966 1180
rect 6092 1027 6158 1180
rect 6284 1027 6350 1180
rect 6476 1027 6542 1180
rect 6668 1027 6734 1180
rect 6860 1027 6926 1180
rect 7344 1027 7410 1180
rect 7536 1027 7602 1180
rect 7728 1027 7794 1180
rect 7920 1027 7986 1180
rect 8112 1027 8178 1180
rect 8304 1027 8370 1180
rect 8496 1027 8562 1180
rect 8688 1027 8754 1180
rect 9172 1027 9238 1180
rect 9364 1027 9430 1180
rect 9556 1027 9622 1180
rect 9748 1027 9814 1180
rect 9940 1027 10006 1180
rect 10132 1027 10198 1180
rect 10324 1027 10390 1180
rect 10516 1027 10582 1180
rect 11000 1027 11066 1180
rect 11192 1027 11258 1180
rect 11384 1027 11450 1180
rect 11576 1027 11642 1180
rect 11768 1027 11834 1180
rect 11960 1027 12026 1180
rect 12152 1027 12218 1180
rect 12344 1027 12410 1180
rect 12828 1027 12894 1180
rect 13020 1027 13086 1180
rect 13212 1027 13278 1180
rect 13404 1027 13470 1180
rect 13596 1027 13662 1180
rect 13788 1027 13854 1180
rect 13980 1027 14046 1180
rect 14172 1027 14238 1180
rect 14656 1027 14722 1180
rect 14848 1027 14914 1180
rect 15040 1027 15106 1180
rect 15232 1027 15298 1180
rect 15424 1027 15490 1180
rect 15616 1027 15682 1180
rect 15808 1027 15874 1180
rect 16000 1027 16066 1180
rect 16484 1027 16550 1180
rect 16676 1027 16742 1180
rect 16868 1027 16934 1180
rect 17060 1027 17126 1180
rect 17252 1027 17318 1180
rect 17444 1027 17510 1180
rect 17636 1027 17702 1180
rect 17828 1027 17894 1180
rect 18312 1027 18378 1180
rect 18504 1027 18570 1180
rect 18696 1027 18762 1180
rect 18888 1027 18954 1180
rect 19080 1027 19146 1180
rect 19272 1027 19338 1180
rect 19464 1027 19530 1180
rect 19656 1027 19722 1180
rect 20140 1027 20206 1180
rect 20332 1027 20398 1180
rect 20524 1027 20590 1180
rect 20716 1027 20782 1180
rect 20908 1027 20974 1180
rect 21100 1027 21166 1180
rect 21292 1027 21358 1180
rect 21484 1027 21550 1180
rect 128 814 194 967
rect 320 814 386 967
rect 512 814 578 967
rect 704 814 770 967
rect 896 814 962 967
rect 1088 814 1154 967
rect 1280 814 1346 967
rect 1472 814 1528 967
rect 1956 814 2022 967
rect 2148 814 2214 967
rect 2340 814 2406 967
rect 2532 814 2598 967
rect 2724 814 2790 967
rect 2916 814 2982 967
rect 3108 814 3174 967
rect 3300 814 3356 967
rect 3784 814 3850 967
rect 3976 814 4042 967
rect 4168 814 4234 967
rect 4360 814 4426 967
rect 4552 814 4618 967
rect 4744 814 4810 967
rect 4936 814 5002 967
rect 5128 814 5184 967
rect 5612 814 5678 967
rect 5804 814 5870 967
rect 5996 814 6062 967
rect 6188 814 6254 967
rect 6380 814 6446 967
rect 6572 814 6638 967
rect 6764 814 6830 967
rect 6956 814 7012 967
rect 7440 814 7506 967
rect 7632 814 7698 967
rect 7824 814 7890 967
rect 8016 814 8082 967
rect 8208 814 8274 967
rect 8400 814 8466 967
rect 8592 814 8658 967
rect 8784 814 8840 967
rect 9268 814 9334 967
rect 9460 814 9526 967
rect 9652 814 9718 967
rect 9844 814 9910 967
rect 10036 814 10102 967
rect 10228 814 10294 967
rect 10420 814 10486 967
rect 10612 814 10668 967
rect 11096 814 11162 967
rect 11288 814 11354 967
rect 11480 814 11546 967
rect 11672 814 11738 967
rect 11864 814 11930 967
rect 12056 814 12122 967
rect 12248 814 12314 967
rect 12440 814 12496 967
rect 12924 814 12990 967
rect 13116 814 13182 967
rect 13308 814 13374 967
rect 13500 814 13566 967
rect 13692 814 13758 967
rect 13884 814 13950 967
rect 14076 814 14142 967
rect 14268 814 14324 967
rect 14752 814 14818 967
rect 14944 814 15010 967
rect 15136 814 15202 967
rect 15328 814 15394 967
rect 15520 814 15586 967
rect 15712 814 15778 967
rect 15904 814 15970 967
rect 16096 814 16152 967
rect 16580 814 16646 967
rect 16772 814 16838 967
rect 16964 814 17030 967
rect 17156 814 17222 967
rect 17348 814 17414 967
rect 17540 814 17606 967
rect 17732 814 17798 967
rect 17924 814 17980 967
rect 18408 814 18474 967
rect 18600 814 18666 967
rect 18792 814 18858 967
rect 18984 814 19050 967
rect 19176 814 19242 967
rect 19368 814 19434 967
rect 19560 814 19626 967
rect 19752 814 19808 967
rect 20236 814 20302 967
rect 20428 814 20494 967
rect 20620 814 20686 967
rect 20812 814 20878 967
rect 21004 814 21070 967
rect 21196 814 21262 967
rect 21388 814 21454 967
rect 21580 814 21636 967
rect 32 313 98 466
rect 224 313 290 466
rect 416 313 482 466
rect 608 313 674 466
rect 800 313 866 466
rect 992 313 1058 466
rect 1184 313 1250 466
rect 1376 313 1442 466
rect 1860 313 1926 466
rect 2052 313 2118 466
rect 2244 313 2310 466
rect 2436 313 2502 466
rect 2628 313 2694 466
rect 2820 313 2886 466
rect 3012 313 3078 466
rect 3204 313 3270 466
rect 3688 313 3754 466
rect 3880 313 3946 466
rect 4072 313 4138 466
rect 4264 313 4330 466
rect 4456 313 4522 466
rect 4648 313 4714 466
rect 4840 313 4906 466
rect 5032 313 5098 466
rect 5516 313 5582 466
rect 5708 313 5774 466
rect 5900 313 5966 466
rect 6092 313 6158 466
rect 6284 313 6350 466
rect 6476 313 6542 466
rect 6668 313 6734 466
rect 6860 313 6926 466
rect 7344 313 7410 466
rect 7536 313 7602 466
rect 7728 313 7794 466
rect 7920 313 7986 466
rect 8112 313 8178 466
rect 8304 313 8370 466
rect 8496 313 8562 466
rect 8688 313 8754 466
rect 9172 313 9238 466
rect 9364 313 9430 466
rect 9556 313 9622 466
rect 9748 313 9814 466
rect 9940 313 10006 466
rect 10132 313 10198 466
rect 10324 313 10390 466
rect 10516 313 10582 466
rect 11000 313 11066 466
rect 11192 313 11258 466
rect 11384 313 11450 466
rect 11576 313 11642 466
rect 11768 313 11834 466
rect 11960 313 12026 466
rect 12152 313 12218 466
rect 12344 313 12410 466
rect 12828 313 12894 466
rect 13020 313 13086 466
rect 13212 313 13278 466
rect 13404 313 13470 466
rect 13596 313 13662 466
rect 13788 313 13854 466
rect 13980 313 14046 466
rect 14172 313 14238 466
rect 14656 313 14722 466
rect 14848 313 14914 466
rect 15040 313 15106 466
rect 15232 313 15298 466
rect 15424 313 15490 466
rect 15616 313 15682 466
rect 15808 313 15874 466
rect 16000 313 16066 466
rect 16484 313 16550 466
rect 16676 313 16742 466
rect 16868 313 16934 466
rect 17060 313 17126 466
rect 17252 313 17318 466
rect 17444 313 17510 466
rect 17636 313 17702 466
rect 17828 313 17894 466
rect 18312 313 18378 466
rect 18504 313 18570 466
rect 18696 313 18762 466
rect 18888 313 18954 466
rect 19080 313 19146 466
rect 19272 313 19338 466
rect 19464 313 19530 466
rect 19656 313 19722 466
rect 20140 313 20206 466
rect 20332 313 20398 466
rect 20524 313 20590 466
rect 20716 313 20782 466
rect 20908 313 20974 466
rect 21100 313 21166 466
rect 21292 313 21358 466
rect 21484 313 21550 466
rect 128 100 194 253
rect 320 100 386 253
rect 512 100 578 253
rect 704 100 770 253
rect 896 100 962 253
rect 1088 100 1154 253
rect 1280 100 1346 253
rect 1472 100 1528 253
rect 1956 100 2022 253
rect 2148 100 2214 253
rect 2340 100 2406 253
rect 2532 100 2598 253
rect 2724 100 2790 253
rect 2916 100 2982 253
rect 3108 100 3174 253
rect 3300 100 3356 253
rect 3784 100 3850 253
rect 3976 100 4042 253
rect 4168 100 4234 253
rect 4360 100 4426 253
rect 4552 100 4618 253
rect 4744 100 4810 253
rect 4936 100 5002 253
rect 5128 100 5184 253
rect 5612 100 5678 253
rect 5804 100 5870 253
rect 5996 100 6062 253
rect 6188 100 6254 253
rect 6380 100 6446 253
rect 6572 100 6638 253
rect 6764 100 6830 253
rect 6956 100 7012 253
rect 7440 100 7506 253
rect 7632 100 7698 253
rect 7824 100 7890 253
rect 8016 100 8082 253
rect 8208 100 8274 253
rect 8400 100 8466 253
rect 8592 100 8658 253
rect 8784 100 8840 253
rect 9268 100 9334 253
rect 9460 100 9526 253
rect 9652 100 9718 253
rect 9844 100 9910 253
rect 10036 100 10102 253
rect 10228 100 10294 253
rect 10420 100 10486 253
rect 10612 100 10668 253
rect 11096 100 11162 253
rect 11288 100 11354 253
rect 11480 100 11546 253
rect 11672 100 11738 253
rect 11864 100 11930 253
rect 12056 100 12122 253
rect 12248 100 12314 253
rect 12440 100 12496 253
rect 12924 100 12990 253
rect 13116 100 13182 253
rect 13308 100 13374 253
rect 13500 100 13566 253
rect 13692 100 13758 253
rect 13884 100 13950 253
rect 14076 100 14142 253
rect 14268 100 14324 253
rect 14752 100 14818 253
rect 14944 100 15010 253
rect 15136 100 15202 253
rect 15328 100 15394 253
rect 15520 100 15586 253
rect 15712 100 15778 253
rect 15904 100 15970 253
rect 16096 100 16152 253
rect 16580 100 16646 253
rect 16772 100 16838 253
rect 16964 100 17030 253
rect 17156 100 17222 253
rect 17348 100 17414 253
rect 17540 100 17606 253
rect 17732 100 17798 253
rect 17924 100 17980 253
rect 18408 100 18474 253
rect 18600 100 18666 253
rect 18792 100 18858 253
rect 18984 100 19050 253
rect 19176 100 19242 253
rect 19368 100 19434 253
rect 19560 100 19626 253
rect 19752 100 19808 253
rect 20236 100 20302 253
rect 20428 100 20494 253
rect 20620 100 20686 253
rect 20812 100 20878 253
rect 21004 100 21070 253
rect 21196 100 21262 253
rect 21388 100 21454 253
rect 21580 100 21636 253
<< metal2 >>
rect 32 21172 98 21182
rect 224 21172 290 21182
rect 416 21172 482 21182
rect 608 21172 674 21182
rect 800 21172 866 21182
rect 992 21172 1058 21182
rect 1184 21172 1250 21182
rect 1376 21172 1442 21182
rect 1860 21172 1926 21182
rect 2052 21172 2118 21182
rect 2244 21172 2310 21182
rect 2436 21172 2502 21182
rect 2628 21172 2694 21182
rect 2820 21172 2886 21182
rect 3012 21172 3078 21182
rect 3204 21172 3270 21182
rect 3688 21172 3754 21182
rect 3880 21172 3946 21182
rect 4072 21172 4138 21182
rect 4264 21172 4330 21182
rect 4456 21172 4522 21182
rect 4648 21172 4714 21182
rect 4840 21172 4906 21182
rect 5032 21172 5098 21182
rect 5516 21172 5582 21182
rect 5708 21172 5774 21182
rect 5900 21172 5966 21182
rect 6092 21172 6158 21182
rect 6284 21172 6350 21182
rect 6476 21172 6542 21182
rect 6668 21172 6734 21182
rect 6860 21172 6926 21182
rect 7344 21172 7410 21182
rect 7536 21172 7602 21182
rect 7728 21172 7794 21182
rect 7920 21172 7986 21182
rect 8112 21172 8178 21182
rect 8304 21172 8370 21182
rect 8496 21172 8562 21182
rect 8688 21172 8754 21182
rect 9172 21172 9238 21182
rect 9364 21172 9430 21182
rect 9556 21172 9622 21182
rect 9748 21172 9814 21182
rect 9940 21172 10006 21182
rect 10132 21172 10198 21182
rect 10324 21172 10390 21182
rect 10516 21172 10582 21182
rect 11000 21172 11066 21182
rect 11192 21172 11258 21182
rect 11384 21172 11450 21182
rect 11576 21172 11642 21182
rect 11768 21172 11834 21182
rect 11960 21172 12026 21182
rect 12152 21172 12218 21182
rect 12344 21172 12410 21182
rect 12828 21172 12894 21182
rect 13020 21172 13086 21182
rect 13212 21172 13278 21182
rect 13404 21172 13470 21182
rect 13596 21172 13662 21182
rect 13788 21172 13854 21182
rect 13980 21172 14046 21182
rect 14172 21172 14238 21182
rect 14656 21172 14722 21182
rect 14848 21172 14914 21182
rect 15040 21172 15106 21182
rect 15232 21172 15298 21182
rect 15424 21172 15490 21182
rect 15616 21172 15682 21182
rect 15808 21172 15874 21182
rect 16000 21172 16066 21182
rect 16484 21172 16550 21182
rect 16676 21172 16742 21182
rect 16868 21172 16934 21182
rect 17060 21172 17126 21182
rect 17252 21172 17318 21182
rect 17444 21172 17510 21182
rect 17636 21172 17702 21182
rect 17828 21172 17894 21182
rect 18312 21172 18378 21182
rect 18504 21172 18570 21182
rect 18696 21172 18762 21182
rect 18888 21172 18954 21182
rect 19080 21172 19146 21182
rect 19272 21172 19338 21182
rect 19464 21172 19530 21182
rect 19656 21172 19722 21182
rect 20140 21172 20206 21182
rect 20332 21172 20398 21182
rect 20524 21172 20590 21182
rect 20716 21172 20782 21182
rect 20908 21172 20974 21182
rect 21100 21172 21166 21182
rect 21292 21172 21358 21182
rect 21484 21172 21550 21182
rect 0 21019 32 21172
rect 98 21019 224 21172
rect 290 21019 416 21172
rect 482 21019 608 21172
rect 674 21019 800 21172
rect 866 21019 992 21172
rect 1058 21019 1184 21172
rect 1250 21019 1376 21172
rect 1828 21019 1860 21172
rect 1926 21019 2052 21172
rect 2118 21019 2244 21172
rect 2310 21019 2436 21172
rect 2502 21019 2628 21172
rect 2694 21019 2820 21172
rect 2886 21019 3012 21172
rect 3078 21019 3204 21172
rect 3656 21019 3688 21172
rect 3754 21019 3880 21172
rect 3946 21019 4072 21172
rect 4138 21019 4264 21172
rect 4330 21019 4456 21172
rect 4522 21019 4648 21172
rect 4714 21019 4840 21172
rect 4906 21019 5032 21172
rect 5484 21019 5516 21172
rect 5582 21019 5708 21172
rect 5774 21019 5900 21172
rect 5966 21019 6092 21172
rect 6158 21019 6284 21172
rect 6350 21019 6476 21172
rect 6542 21019 6668 21172
rect 6734 21019 6860 21172
rect 7312 21019 7344 21172
rect 7410 21019 7536 21172
rect 7602 21019 7728 21172
rect 7794 21019 7920 21172
rect 7986 21019 8112 21172
rect 8178 21019 8304 21172
rect 8370 21019 8496 21172
rect 8562 21019 8688 21172
rect 9140 21019 9172 21172
rect 9238 21019 9364 21172
rect 9430 21019 9556 21172
rect 9622 21019 9748 21172
rect 9814 21019 9940 21172
rect 10006 21019 10132 21172
rect 10198 21019 10324 21172
rect 10390 21019 10516 21172
rect 10968 21019 11000 21172
rect 11066 21019 11192 21172
rect 11258 21019 11384 21172
rect 11450 21019 11576 21172
rect 11642 21019 11768 21172
rect 11834 21019 11960 21172
rect 12026 21019 12152 21172
rect 12218 21019 12344 21172
rect 12796 21019 12828 21172
rect 12894 21019 13020 21172
rect 13086 21019 13212 21172
rect 13278 21019 13404 21172
rect 13470 21019 13596 21172
rect 13662 21019 13788 21172
rect 13854 21019 13980 21172
rect 14046 21019 14172 21172
rect 14624 21019 14656 21172
rect 14722 21019 14848 21172
rect 14914 21019 15040 21172
rect 15106 21019 15232 21172
rect 15298 21019 15424 21172
rect 15490 21019 15616 21172
rect 15682 21019 15808 21172
rect 15874 21019 16000 21172
rect 16452 21019 16484 21172
rect 16550 21019 16676 21172
rect 16742 21019 16868 21172
rect 16934 21019 17060 21172
rect 17126 21019 17252 21172
rect 17318 21019 17444 21172
rect 17510 21019 17636 21172
rect 17702 21019 17828 21172
rect 18280 21019 18312 21172
rect 18378 21019 18504 21172
rect 18570 21019 18696 21172
rect 18762 21019 18888 21172
rect 18954 21019 19080 21172
rect 19146 21019 19272 21172
rect 19338 21019 19464 21172
rect 19530 21019 19656 21172
rect 20108 21019 20140 21172
rect 20206 21019 20332 21172
rect 20398 21019 20524 21172
rect 20590 21019 20716 21172
rect 20782 21019 20908 21172
rect 20974 21019 21100 21172
rect 21166 21019 21292 21172
rect 21358 21019 21484 21172
rect 32 21009 98 21019
rect 224 21009 290 21019
rect 416 21009 482 21019
rect 608 21009 674 21019
rect 800 21009 866 21019
rect 992 21009 1058 21019
rect 1184 21009 1250 21019
rect 1376 21009 1442 21019
rect 1860 21009 1926 21019
rect 2052 21009 2118 21019
rect 2244 21009 2310 21019
rect 2436 21009 2502 21019
rect 2628 21009 2694 21019
rect 2820 21009 2886 21019
rect 3012 21009 3078 21019
rect 3204 21009 3270 21019
rect 3688 21009 3754 21019
rect 3880 21009 3946 21019
rect 4072 21009 4138 21019
rect 4264 21009 4330 21019
rect 4456 21009 4522 21019
rect 4648 21009 4714 21019
rect 4840 21009 4906 21019
rect 5032 21009 5098 21019
rect 5516 21009 5582 21019
rect 5708 21009 5774 21019
rect 5900 21009 5966 21019
rect 6092 21009 6158 21019
rect 6284 21009 6350 21019
rect 6476 21009 6542 21019
rect 6668 21009 6734 21019
rect 6860 21009 6926 21019
rect 7344 21009 7410 21019
rect 7536 21009 7602 21019
rect 7728 21009 7794 21019
rect 7920 21009 7986 21019
rect 8112 21009 8178 21019
rect 8304 21009 8370 21019
rect 8496 21009 8562 21019
rect 8688 21009 8754 21019
rect 9172 21009 9238 21019
rect 9364 21009 9430 21019
rect 9556 21009 9622 21019
rect 9748 21009 9814 21019
rect 9940 21009 10006 21019
rect 10132 21009 10198 21019
rect 10324 21009 10390 21019
rect 10516 21009 10582 21019
rect 11000 21009 11066 21019
rect 11192 21009 11258 21019
rect 11384 21009 11450 21019
rect 11576 21009 11642 21019
rect 11768 21009 11834 21019
rect 11960 21009 12026 21019
rect 12152 21009 12218 21019
rect 12344 21009 12410 21019
rect 12828 21009 12894 21019
rect 13020 21009 13086 21019
rect 13212 21009 13278 21019
rect 13404 21009 13470 21019
rect 13596 21009 13662 21019
rect 13788 21009 13854 21019
rect 13980 21009 14046 21019
rect 14172 21009 14238 21019
rect 14656 21009 14722 21019
rect 14848 21009 14914 21019
rect 15040 21009 15106 21019
rect 15232 21009 15298 21019
rect 15424 21009 15490 21019
rect 15616 21009 15682 21019
rect 15808 21009 15874 21019
rect 16000 21009 16066 21019
rect 16484 21009 16550 21019
rect 16676 21009 16742 21019
rect 16868 21009 16934 21019
rect 17060 21009 17126 21019
rect 17252 21009 17318 21019
rect 17444 21009 17510 21019
rect 17636 21009 17702 21019
rect 17828 21009 17894 21019
rect 18312 21009 18378 21019
rect 18504 21009 18570 21019
rect 18696 21009 18762 21019
rect 18888 21009 18954 21019
rect 19080 21009 19146 21019
rect 19272 21009 19338 21019
rect 19464 21009 19530 21019
rect 19656 21009 19722 21019
rect 20140 21009 20206 21019
rect 20332 21009 20398 21019
rect 20524 21009 20590 21019
rect 20716 21009 20782 21019
rect 20908 21009 20974 21019
rect 21100 21009 21166 21019
rect 21292 21009 21358 21019
rect 21484 21009 21550 21019
rect 128 20959 194 20969
rect 320 20959 386 20969
rect 512 20959 578 20969
rect 704 20959 770 20969
rect 896 20959 962 20969
rect 1088 20959 1154 20969
rect 1280 20959 1346 20969
rect 1472 20959 1528 20969
rect 1956 20959 2022 20969
rect 2148 20959 2214 20969
rect 2340 20959 2406 20969
rect 2532 20959 2598 20969
rect 2724 20959 2790 20969
rect 2916 20959 2982 20969
rect 3108 20959 3174 20969
rect 3300 20959 3356 20969
rect 3784 20959 3850 20969
rect 3976 20959 4042 20969
rect 4168 20959 4234 20969
rect 4360 20959 4426 20969
rect 4552 20959 4618 20969
rect 4744 20959 4810 20969
rect 4936 20959 5002 20969
rect 5128 20959 5184 20969
rect 5612 20959 5678 20969
rect 5804 20959 5870 20969
rect 5996 20959 6062 20969
rect 6188 20959 6254 20969
rect 6380 20959 6446 20969
rect 6572 20959 6638 20969
rect 6764 20959 6830 20969
rect 6956 20959 7012 20969
rect 7440 20959 7506 20969
rect 7632 20959 7698 20969
rect 7824 20959 7890 20969
rect 8016 20959 8082 20969
rect 8208 20959 8274 20969
rect 8400 20959 8466 20969
rect 8592 20959 8658 20969
rect 8784 20959 8840 20969
rect 9268 20959 9334 20969
rect 9460 20959 9526 20969
rect 9652 20959 9718 20969
rect 9844 20959 9910 20969
rect 10036 20959 10102 20969
rect 10228 20959 10294 20969
rect 10420 20959 10486 20969
rect 10612 20959 10668 20969
rect 11096 20959 11162 20969
rect 11288 20959 11354 20969
rect 11480 20959 11546 20969
rect 11672 20959 11738 20969
rect 11864 20959 11930 20969
rect 12056 20959 12122 20969
rect 12248 20959 12314 20969
rect 12440 20959 12496 20969
rect 12924 20959 12990 20969
rect 13116 20959 13182 20969
rect 13308 20959 13374 20969
rect 13500 20959 13566 20969
rect 13692 20959 13758 20969
rect 13884 20959 13950 20969
rect 14076 20959 14142 20969
rect 14268 20959 14324 20969
rect 14752 20959 14818 20969
rect 14944 20959 15010 20969
rect 15136 20959 15202 20969
rect 15328 20959 15394 20969
rect 15520 20959 15586 20969
rect 15712 20959 15778 20969
rect 15904 20959 15970 20969
rect 16096 20959 16152 20969
rect 16580 20959 16646 20969
rect 16772 20959 16838 20969
rect 16964 20959 17030 20969
rect 17156 20959 17222 20969
rect 17348 20959 17414 20969
rect 17540 20959 17606 20969
rect 17732 20959 17798 20969
rect 17924 20959 17980 20969
rect 18408 20959 18474 20969
rect 18600 20959 18666 20969
rect 18792 20959 18858 20969
rect 18984 20959 19050 20969
rect 19176 20959 19242 20969
rect 19368 20959 19434 20969
rect 19560 20959 19626 20969
rect 19752 20959 19808 20969
rect 20236 20959 20302 20969
rect 20428 20959 20494 20969
rect 20620 20959 20686 20969
rect 20812 20959 20878 20969
rect 21004 20959 21070 20969
rect 21196 20959 21262 20969
rect 21388 20959 21454 20969
rect 21580 20959 21636 20969
rect 0 20806 128 20959
rect 194 20806 320 20959
rect 386 20806 512 20959
rect 578 20806 704 20959
rect 770 20806 896 20959
rect 962 20806 1088 20959
rect 1154 20806 1280 20959
rect 1346 20806 1472 20959
rect 1528 20806 1708 20959
rect 1828 20806 1956 20959
rect 2022 20806 2148 20959
rect 2214 20806 2340 20959
rect 2406 20806 2532 20959
rect 2598 20806 2724 20959
rect 2790 20806 2916 20959
rect 2982 20806 3108 20959
rect 3174 20806 3300 20959
rect 3356 20806 3536 20959
rect 3656 20806 3784 20959
rect 3850 20806 3976 20959
rect 4042 20806 4168 20959
rect 4234 20806 4360 20959
rect 4426 20806 4552 20959
rect 4618 20806 4744 20959
rect 4810 20806 4936 20959
rect 5002 20806 5128 20959
rect 5184 20806 5364 20959
rect 5484 20806 5612 20959
rect 5678 20806 5804 20959
rect 5870 20806 5996 20959
rect 6062 20806 6188 20959
rect 6254 20806 6380 20959
rect 6446 20806 6572 20959
rect 6638 20806 6764 20959
rect 6830 20806 6956 20959
rect 7012 20806 7192 20959
rect 7312 20806 7440 20959
rect 7506 20806 7632 20959
rect 7698 20806 7824 20959
rect 7890 20806 8016 20959
rect 8082 20806 8208 20959
rect 8274 20806 8400 20959
rect 8466 20806 8592 20959
rect 8658 20806 8784 20959
rect 8840 20806 9020 20959
rect 9140 20806 9268 20959
rect 9334 20806 9460 20959
rect 9526 20806 9652 20959
rect 9718 20806 9844 20959
rect 9910 20806 10036 20959
rect 10102 20806 10228 20959
rect 10294 20806 10420 20959
rect 10486 20806 10612 20959
rect 10668 20806 10848 20959
rect 10968 20806 11096 20959
rect 11162 20806 11288 20959
rect 11354 20806 11480 20959
rect 11546 20806 11672 20959
rect 11738 20806 11864 20959
rect 11930 20806 12056 20959
rect 12122 20806 12248 20959
rect 12314 20806 12440 20959
rect 12496 20806 12676 20959
rect 12796 20806 12924 20959
rect 12990 20806 13116 20959
rect 13182 20806 13308 20959
rect 13374 20806 13500 20959
rect 13566 20806 13692 20959
rect 13758 20806 13884 20959
rect 13950 20806 14076 20959
rect 14142 20806 14268 20959
rect 14324 20806 14504 20959
rect 14624 20806 14752 20959
rect 14818 20806 14944 20959
rect 15010 20806 15136 20959
rect 15202 20806 15328 20959
rect 15394 20806 15520 20959
rect 15586 20806 15712 20959
rect 15778 20806 15904 20959
rect 15970 20806 16096 20959
rect 16152 20806 16332 20959
rect 16452 20806 16580 20959
rect 16646 20806 16772 20959
rect 16838 20806 16964 20959
rect 17030 20806 17156 20959
rect 17222 20806 17348 20959
rect 17414 20806 17540 20959
rect 17606 20806 17732 20959
rect 17798 20806 17924 20959
rect 17980 20806 18160 20959
rect 18280 20806 18408 20959
rect 18474 20806 18600 20959
rect 18666 20806 18792 20959
rect 18858 20806 18984 20959
rect 19050 20806 19176 20959
rect 19242 20806 19368 20959
rect 19434 20806 19560 20959
rect 19626 20806 19752 20959
rect 19808 20806 19988 20959
rect 20108 20806 20236 20959
rect 20302 20806 20428 20959
rect 20494 20806 20620 20959
rect 20686 20806 20812 20959
rect 20878 20806 21004 20959
rect 21070 20806 21196 20959
rect 21262 20806 21388 20959
rect 21454 20806 21580 20959
rect 21636 20806 21816 20959
rect 128 20796 194 20806
rect 320 20796 386 20806
rect 512 20796 578 20806
rect 704 20796 770 20806
rect 896 20796 962 20806
rect 1088 20796 1154 20806
rect 1280 20796 1346 20806
rect 1472 20796 1528 20806
rect 1956 20796 2022 20806
rect 2148 20796 2214 20806
rect 2340 20796 2406 20806
rect 2532 20796 2598 20806
rect 2724 20796 2790 20806
rect 2916 20796 2982 20806
rect 3108 20796 3174 20806
rect 3300 20796 3356 20806
rect 3784 20796 3850 20806
rect 3976 20796 4042 20806
rect 4168 20796 4234 20806
rect 4360 20796 4426 20806
rect 4552 20796 4618 20806
rect 4744 20796 4810 20806
rect 4936 20796 5002 20806
rect 5128 20796 5184 20806
rect 5612 20796 5678 20806
rect 5804 20796 5870 20806
rect 5996 20796 6062 20806
rect 6188 20796 6254 20806
rect 6380 20796 6446 20806
rect 6572 20796 6638 20806
rect 6764 20796 6830 20806
rect 6956 20796 7012 20806
rect 7440 20796 7506 20806
rect 7632 20796 7698 20806
rect 7824 20796 7890 20806
rect 8016 20796 8082 20806
rect 8208 20796 8274 20806
rect 8400 20796 8466 20806
rect 8592 20796 8658 20806
rect 8784 20796 8840 20806
rect 9268 20796 9334 20806
rect 9460 20796 9526 20806
rect 9652 20796 9718 20806
rect 9844 20796 9910 20806
rect 10036 20796 10102 20806
rect 10228 20796 10294 20806
rect 10420 20796 10486 20806
rect 10612 20796 10668 20806
rect 11096 20796 11162 20806
rect 11288 20796 11354 20806
rect 11480 20796 11546 20806
rect 11672 20796 11738 20806
rect 11864 20796 11930 20806
rect 12056 20796 12122 20806
rect 12248 20796 12314 20806
rect 12440 20796 12496 20806
rect 12924 20796 12990 20806
rect 13116 20796 13182 20806
rect 13308 20796 13374 20806
rect 13500 20796 13566 20806
rect 13692 20796 13758 20806
rect 13884 20796 13950 20806
rect 14076 20796 14142 20806
rect 14268 20796 14324 20806
rect 14752 20796 14818 20806
rect 14944 20796 15010 20806
rect 15136 20796 15202 20806
rect 15328 20796 15394 20806
rect 15520 20796 15586 20806
rect 15712 20796 15778 20806
rect 15904 20796 15970 20806
rect 16096 20796 16152 20806
rect 16580 20796 16646 20806
rect 16772 20796 16838 20806
rect 16964 20796 17030 20806
rect 17156 20796 17222 20806
rect 17348 20796 17414 20806
rect 17540 20796 17606 20806
rect 17732 20796 17798 20806
rect 17924 20796 17980 20806
rect 18408 20796 18474 20806
rect 18600 20796 18666 20806
rect 18792 20796 18858 20806
rect 18984 20796 19050 20806
rect 19176 20796 19242 20806
rect 19368 20796 19434 20806
rect 19560 20796 19626 20806
rect 19752 20796 19808 20806
rect 20236 20796 20302 20806
rect 20428 20796 20494 20806
rect 20620 20796 20686 20806
rect 20812 20796 20878 20806
rect 21004 20796 21070 20806
rect 21196 20796 21262 20806
rect 21388 20796 21454 20806
rect 21580 20796 21636 20806
rect 32 20458 98 20468
rect 224 20458 290 20468
rect 416 20458 482 20468
rect 608 20458 674 20468
rect 800 20458 866 20468
rect 992 20458 1058 20468
rect 1184 20458 1250 20468
rect 1376 20458 1442 20468
rect 1860 20458 1926 20468
rect 2052 20458 2118 20468
rect 2244 20458 2310 20468
rect 2436 20458 2502 20468
rect 2628 20458 2694 20468
rect 2820 20458 2886 20468
rect 3012 20458 3078 20468
rect 3204 20458 3270 20468
rect 3688 20458 3754 20468
rect 3880 20458 3946 20468
rect 4072 20458 4138 20468
rect 4264 20458 4330 20468
rect 4456 20458 4522 20468
rect 4648 20458 4714 20468
rect 4840 20458 4906 20468
rect 5032 20458 5098 20468
rect 5516 20458 5582 20468
rect 5708 20458 5774 20468
rect 5900 20458 5966 20468
rect 6092 20458 6158 20468
rect 6284 20458 6350 20468
rect 6476 20458 6542 20468
rect 6668 20458 6734 20468
rect 6860 20458 6926 20468
rect 7344 20458 7410 20468
rect 7536 20458 7602 20468
rect 7728 20458 7794 20468
rect 7920 20458 7986 20468
rect 8112 20458 8178 20468
rect 8304 20458 8370 20468
rect 8496 20458 8562 20468
rect 8688 20458 8754 20468
rect 9172 20458 9238 20468
rect 9364 20458 9430 20468
rect 9556 20458 9622 20468
rect 9748 20458 9814 20468
rect 9940 20458 10006 20468
rect 10132 20458 10198 20468
rect 10324 20458 10390 20468
rect 10516 20458 10582 20468
rect 11000 20458 11066 20468
rect 11192 20458 11258 20468
rect 11384 20458 11450 20468
rect 11576 20458 11642 20468
rect 11768 20458 11834 20468
rect 11960 20458 12026 20468
rect 12152 20458 12218 20468
rect 12344 20458 12410 20468
rect 12828 20458 12894 20468
rect 13020 20458 13086 20468
rect 13212 20458 13278 20468
rect 13404 20458 13470 20468
rect 13596 20458 13662 20468
rect 13788 20458 13854 20468
rect 13980 20458 14046 20468
rect 14172 20458 14238 20468
rect 14656 20458 14722 20468
rect 14848 20458 14914 20468
rect 15040 20458 15106 20468
rect 15232 20458 15298 20468
rect 15424 20458 15490 20468
rect 15616 20458 15682 20468
rect 15808 20458 15874 20468
rect 16000 20458 16066 20468
rect 16484 20458 16550 20468
rect 16676 20458 16742 20468
rect 16868 20458 16934 20468
rect 17060 20458 17126 20468
rect 17252 20458 17318 20468
rect 17444 20458 17510 20468
rect 17636 20458 17702 20468
rect 17828 20458 17894 20468
rect 18312 20458 18378 20468
rect 18504 20458 18570 20468
rect 18696 20458 18762 20468
rect 18888 20458 18954 20468
rect 19080 20458 19146 20468
rect 19272 20458 19338 20468
rect 19464 20458 19530 20468
rect 19656 20458 19722 20468
rect 20140 20458 20206 20468
rect 20332 20458 20398 20468
rect 20524 20458 20590 20468
rect 20716 20458 20782 20468
rect 20908 20458 20974 20468
rect 21100 20458 21166 20468
rect 21292 20458 21358 20468
rect 21484 20458 21550 20468
rect 0 20305 32 20458
rect 98 20305 224 20458
rect 290 20305 416 20458
rect 482 20305 608 20458
rect 674 20305 800 20458
rect 866 20305 992 20458
rect 1058 20305 1184 20458
rect 1250 20305 1376 20458
rect 1828 20305 1860 20458
rect 1926 20305 2052 20458
rect 2118 20305 2244 20458
rect 2310 20305 2436 20458
rect 2502 20305 2628 20458
rect 2694 20305 2820 20458
rect 2886 20305 3012 20458
rect 3078 20305 3204 20458
rect 3656 20305 3688 20458
rect 3754 20305 3880 20458
rect 3946 20305 4072 20458
rect 4138 20305 4264 20458
rect 4330 20305 4456 20458
rect 4522 20305 4648 20458
rect 4714 20305 4840 20458
rect 4906 20305 5032 20458
rect 5484 20305 5516 20458
rect 5582 20305 5708 20458
rect 5774 20305 5900 20458
rect 5966 20305 6092 20458
rect 6158 20305 6284 20458
rect 6350 20305 6476 20458
rect 6542 20305 6668 20458
rect 6734 20305 6860 20458
rect 7312 20305 7344 20458
rect 7410 20305 7536 20458
rect 7602 20305 7728 20458
rect 7794 20305 7920 20458
rect 7986 20305 8112 20458
rect 8178 20305 8304 20458
rect 8370 20305 8496 20458
rect 8562 20305 8688 20458
rect 9140 20305 9172 20458
rect 9238 20305 9364 20458
rect 9430 20305 9556 20458
rect 9622 20305 9748 20458
rect 9814 20305 9940 20458
rect 10006 20305 10132 20458
rect 10198 20305 10324 20458
rect 10390 20305 10516 20458
rect 10968 20305 11000 20458
rect 11066 20305 11192 20458
rect 11258 20305 11384 20458
rect 11450 20305 11576 20458
rect 11642 20305 11768 20458
rect 11834 20305 11960 20458
rect 12026 20305 12152 20458
rect 12218 20305 12344 20458
rect 12796 20305 12828 20458
rect 12894 20305 13020 20458
rect 13086 20305 13212 20458
rect 13278 20305 13404 20458
rect 13470 20305 13596 20458
rect 13662 20305 13788 20458
rect 13854 20305 13980 20458
rect 14046 20305 14172 20458
rect 14624 20305 14656 20458
rect 14722 20305 14848 20458
rect 14914 20305 15040 20458
rect 15106 20305 15232 20458
rect 15298 20305 15424 20458
rect 15490 20305 15616 20458
rect 15682 20305 15808 20458
rect 15874 20305 16000 20458
rect 16452 20305 16484 20458
rect 16550 20305 16676 20458
rect 16742 20305 16868 20458
rect 16934 20305 17060 20458
rect 17126 20305 17252 20458
rect 17318 20305 17444 20458
rect 17510 20305 17636 20458
rect 17702 20305 17828 20458
rect 18280 20305 18312 20458
rect 18378 20305 18504 20458
rect 18570 20305 18696 20458
rect 18762 20305 18888 20458
rect 18954 20305 19080 20458
rect 19146 20305 19272 20458
rect 19338 20305 19464 20458
rect 19530 20305 19656 20458
rect 20108 20305 20140 20458
rect 20206 20305 20332 20458
rect 20398 20305 20524 20458
rect 20590 20305 20716 20458
rect 20782 20305 20908 20458
rect 20974 20305 21100 20458
rect 21166 20305 21292 20458
rect 21358 20305 21484 20458
rect 32 20295 98 20305
rect 224 20295 290 20305
rect 416 20295 482 20305
rect 608 20295 674 20305
rect 800 20295 866 20305
rect 992 20295 1058 20305
rect 1184 20295 1250 20305
rect 1376 20295 1442 20305
rect 1860 20295 1926 20305
rect 2052 20295 2118 20305
rect 2244 20295 2310 20305
rect 2436 20295 2502 20305
rect 2628 20295 2694 20305
rect 2820 20295 2886 20305
rect 3012 20295 3078 20305
rect 3204 20295 3270 20305
rect 3688 20295 3754 20305
rect 3880 20295 3946 20305
rect 4072 20295 4138 20305
rect 4264 20295 4330 20305
rect 4456 20295 4522 20305
rect 4648 20295 4714 20305
rect 4840 20295 4906 20305
rect 5032 20295 5098 20305
rect 5516 20295 5582 20305
rect 5708 20295 5774 20305
rect 5900 20295 5966 20305
rect 6092 20295 6158 20305
rect 6284 20295 6350 20305
rect 6476 20295 6542 20305
rect 6668 20295 6734 20305
rect 6860 20295 6926 20305
rect 7344 20295 7410 20305
rect 7536 20295 7602 20305
rect 7728 20295 7794 20305
rect 7920 20295 7986 20305
rect 8112 20295 8178 20305
rect 8304 20295 8370 20305
rect 8496 20295 8562 20305
rect 8688 20295 8754 20305
rect 9172 20295 9238 20305
rect 9364 20295 9430 20305
rect 9556 20295 9622 20305
rect 9748 20295 9814 20305
rect 9940 20295 10006 20305
rect 10132 20295 10198 20305
rect 10324 20295 10390 20305
rect 10516 20295 10582 20305
rect 11000 20295 11066 20305
rect 11192 20295 11258 20305
rect 11384 20295 11450 20305
rect 11576 20295 11642 20305
rect 11768 20295 11834 20305
rect 11960 20295 12026 20305
rect 12152 20295 12218 20305
rect 12344 20295 12410 20305
rect 12828 20295 12894 20305
rect 13020 20295 13086 20305
rect 13212 20295 13278 20305
rect 13404 20295 13470 20305
rect 13596 20295 13662 20305
rect 13788 20295 13854 20305
rect 13980 20295 14046 20305
rect 14172 20295 14238 20305
rect 14656 20295 14722 20305
rect 14848 20295 14914 20305
rect 15040 20295 15106 20305
rect 15232 20295 15298 20305
rect 15424 20295 15490 20305
rect 15616 20295 15682 20305
rect 15808 20295 15874 20305
rect 16000 20295 16066 20305
rect 16484 20295 16550 20305
rect 16676 20295 16742 20305
rect 16868 20295 16934 20305
rect 17060 20295 17126 20305
rect 17252 20295 17318 20305
rect 17444 20295 17510 20305
rect 17636 20295 17702 20305
rect 17828 20295 17894 20305
rect 18312 20295 18378 20305
rect 18504 20295 18570 20305
rect 18696 20295 18762 20305
rect 18888 20295 18954 20305
rect 19080 20295 19146 20305
rect 19272 20295 19338 20305
rect 19464 20295 19530 20305
rect 19656 20295 19722 20305
rect 20140 20295 20206 20305
rect 20332 20295 20398 20305
rect 20524 20295 20590 20305
rect 20716 20295 20782 20305
rect 20908 20295 20974 20305
rect 21100 20295 21166 20305
rect 21292 20295 21358 20305
rect 21484 20295 21550 20305
rect 128 20245 194 20255
rect 320 20245 386 20255
rect 512 20245 578 20255
rect 704 20245 770 20255
rect 896 20245 962 20255
rect 1088 20245 1154 20255
rect 1280 20245 1346 20255
rect 1472 20245 1528 20255
rect 1956 20245 2022 20255
rect 2148 20245 2214 20255
rect 2340 20245 2406 20255
rect 2532 20245 2598 20255
rect 2724 20245 2790 20255
rect 2916 20245 2982 20255
rect 3108 20245 3174 20255
rect 3300 20245 3356 20255
rect 3784 20245 3850 20255
rect 3976 20245 4042 20255
rect 4168 20245 4234 20255
rect 4360 20245 4426 20255
rect 4552 20245 4618 20255
rect 4744 20245 4810 20255
rect 4936 20245 5002 20255
rect 5128 20245 5184 20255
rect 5612 20245 5678 20255
rect 5804 20245 5870 20255
rect 5996 20245 6062 20255
rect 6188 20245 6254 20255
rect 6380 20245 6446 20255
rect 6572 20245 6638 20255
rect 6764 20245 6830 20255
rect 6956 20245 7012 20255
rect 7440 20245 7506 20255
rect 7632 20245 7698 20255
rect 7824 20245 7890 20255
rect 8016 20245 8082 20255
rect 8208 20245 8274 20255
rect 8400 20245 8466 20255
rect 8592 20245 8658 20255
rect 8784 20245 8840 20255
rect 9268 20245 9334 20255
rect 9460 20245 9526 20255
rect 9652 20245 9718 20255
rect 9844 20245 9910 20255
rect 10036 20245 10102 20255
rect 10228 20245 10294 20255
rect 10420 20245 10486 20255
rect 10612 20245 10668 20255
rect 11096 20245 11162 20255
rect 11288 20245 11354 20255
rect 11480 20245 11546 20255
rect 11672 20245 11738 20255
rect 11864 20245 11930 20255
rect 12056 20245 12122 20255
rect 12248 20245 12314 20255
rect 12440 20245 12496 20255
rect 12924 20245 12990 20255
rect 13116 20245 13182 20255
rect 13308 20245 13374 20255
rect 13500 20245 13566 20255
rect 13692 20245 13758 20255
rect 13884 20245 13950 20255
rect 14076 20245 14142 20255
rect 14268 20245 14324 20255
rect 14752 20245 14818 20255
rect 14944 20245 15010 20255
rect 15136 20245 15202 20255
rect 15328 20245 15394 20255
rect 15520 20245 15586 20255
rect 15712 20245 15778 20255
rect 15904 20245 15970 20255
rect 16096 20245 16152 20255
rect 16580 20245 16646 20255
rect 16772 20245 16838 20255
rect 16964 20245 17030 20255
rect 17156 20245 17222 20255
rect 17348 20245 17414 20255
rect 17540 20245 17606 20255
rect 17732 20245 17798 20255
rect 17924 20245 17980 20255
rect 18408 20245 18474 20255
rect 18600 20245 18666 20255
rect 18792 20245 18858 20255
rect 18984 20245 19050 20255
rect 19176 20245 19242 20255
rect 19368 20245 19434 20255
rect 19560 20245 19626 20255
rect 19752 20245 19808 20255
rect 20236 20245 20302 20255
rect 20428 20245 20494 20255
rect 20620 20245 20686 20255
rect 20812 20245 20878 20255
rect 21004 20245 21070 20255
rect 21196 20245 21262 20255
rect 21388 20245 21454 20255
rect 21580 20245 21636 20255
rect 0 20092 128 20245
rect 194 20092 320 20245
rect 386 20092 512 20245
rect 578 20092 704 20245
rect 770 20092 896 20245
rect 962 20092 1088 20245
rect 1154 20092 1280 20245
rect 1346 20092 1472 20245
rect 1528 20092 1708 20245
rect 1828 20092 1956 20245
rect 2022 20092 2148 20245
rect 2214 20092 2340 20245
rect 2406 20092 2532 20245
rect 2598 20092 2724 20245
rect 2790 20092 2916 20245
rect 2982 20092 3108 20245
rect 3174 20092 3300 20245
rect 3356 20092 3536 20245
rect 3656 20092 3784 20245
rect 3850 20092 3976 20245
rect 4042 20092 4168 20245
rect 4234 20092 4360 20245
rect 4426 20092 4552 20245
rect 4618 20092 4744 20245
rect 4810 20092 4936 20245
rect 5002 20092 5128 20245
rect 5184 20092 5364 20245
rect 5484 20092 5612 20245
rect 5678 20092 5804 20245
rect 5870 20092 5996 20245
rect 6062 20092 6188 20245
rect 6254 20092 6380 20245
rect 6446 20092 6572 20245
rect 6638 20092 6764 20245
rect 6830 20092 6956 20245
rect 7012 20092 7192 20245
rect 7312 20092 7440 20245
rect 7506 20092 7632 20245
rect 7698 20092 7824 20245
rect 7890 20092 8016 20245
rect 8082 20092 8208 20245
rect 8274 20092 8400 20245
rect 8466 20092 8592 20245
rect 8658 20092 8784 20245
rect 8840 20092 9020 20245
rect 9140 20092 9268 20245
rect 9334 20092 9460 20245
rect 9526 20092 9652 20245
rect 9718 20092 9844 20245
rect 9910 20092 10036 20245
rect 10102 20092 10228 20245
rect 10294 20092 10420 20245
rect 10486 20092 10612 20245
rect 10668 20092 10848 20245
rect 10968 20092 11096 20245
rect 11162 20092 11288 20245
rect 11354 20092 11480 20245
rect 11546 20092 11672 20245
rect 11738 20092 11864 20245
rect 11930 20092 12056 20245
rect 12122 20092 12248 20245
rect 12314 20092 12440 20245
rect 12496 20092 12676 20245
rect 12796 20092 12924 20245
rect 12990 20092 13116 20245
rect 13182 20092 13308 20245
rect 13374 20092 13500 20245
rect 13566 20092 13692 20245
rect 13758 20092 13884 20245
rect 13950 20092 14076 20245
rect 14142 20092 14268 20245
rect 14324 20092 14504 20245
rect 14624 20092 14752 20245
rect 14818 20092 14944 20245
rect 15010 20092 15136 20245
rect 15202 20092 15328 20245
rect 15394 20092 15520 20245
rect 15586 20092 15712 20245
rect 15778 20092 15904 20245
rect 15970 20092 16096 20245
rect 16152 20092 16332 20245
rect 16452 20092 16580 20245
rect 16646 20092 16772 20245
rect 16838 20092 16964 20245
rect 17030 20092 17156 20245
rect 17222 20092 17348 20245
rect 17414 20092 17540 20245
rect 17606 20092 17732 20245
rect 17798 20092 17924 20245
rect 17980 20092 18160 20245
rect 18280 20092 18408 20245
rect 18474 20092 18600 20245
rect 18666 20092 18792 20245
rect 18858 20092 18984 20245
rect 19050 20092 19176 20245
rect 19242 20092 19368 20245
rect 19434 20092 19560 20245
rect 19626 20092 19752 20245
rect 19808 20092 19988 20245
rect 20108 20092 20236 20245
rect 20302 20092 20428 20245
rect 20494 20092 20620 20245
rect 20686 20092 20812 20245
rect 20878 20092 21004 20245
rect 21070 20092 21196 20245
rect 21262 20092 21388 20245
rect 21454 20092 21580 20245
rect 21636 20092 21816 20245
rect 128 20082 194 20092
rect 320 20082 386 20092
rect 512 20082 578 20092
rect 704 20082 770 20092
rect 896 20082 962 20092
rect 1088 20082 1154 20092
rect 1280 20082 1346 20092
rect 1472 20082 1528 20092
rect 1956 20082 2022 20092
rect 2148 20082 2214 20092
rect 2340 20082 2406 20092
rect 2532 20082 2598 20092
rect 2724 20082 2790 20092
rect 2916 20082 2982 20092
rect 3108 20082 3174 20092
rect 3300 20082 3356 20092
rect 3784 20082 3850 20092
rect 3976 20082 4042 20092
rect 4168 20082 4234 20092
rect 4360 20082 4426 20092
rect 4552 20082 4618 20092
rect 4744 20082 4810 20092
rect 4936 20082 5002 20092
rect 5128 20082 5184 20092
rect 5612 20082 5678 20092
rect 5804 20082 5870 20092
rect 5996 20082 6062 20092
rect 6188 20082 6254 20092
rect 6380 20082 6446 20092
rect 6572 20082 6638 20092
rect 6764 20082 6830 20092
rect 6956 20082 7012 20092
rect 7440 20082 7506 20092
rect 7632 20082 7698 20092
rect 7824 20082 7890 20092
rect 8016 20082 8082 20092
rect 8208 20082 8274 20092
rect 8400 20082 8466 20092
rect 8592 20082 8658 20092
rect 8784 20082 8840 20092
rect 9268 20082 9334 20092
rect 9460 20082 9526 20092
rect 9652 20082 9718 20092
rect 9844 20082 9910 20092
rect 10036 20082 10102 20092
rect 10228 20082 10294 20092
rect 10420 20082 10486 20092
rect 10612 20082 10668 20092
rect 11096 20082 11162 20092
rect 11288 20082 11354 20092
rect 11480 20082 11546 20092
rect 11672 20082 11738 20092
rect 11864 20082 11930 20092
rect 12056 20082 12122 20092
rect 12248 20082 12314 20092
rect 12440 20082 12496 20092
rect 12924 20082 12990 20092
rect 13116 20082 13182 20092
rect 13308 20082 13374 20092
rect 13500 20082 13566 20092
rect 13692 20082 13758 20092
rect 13884 20082 13950 20092
rect 14076 20082 14142 20092
rect 14268 20082 14324 20092
rect 14752 20082 14818 20092
rect 14944 20082 15010 20092
rect 15136 20082 15202 20092
rect 15328 20082 15394 20092
rect 15520 20082 15586 20092
rect 15712 20082 15778 20092
rect 15904 20082 15970 20092
rect 16096 20082 16152 20092
rect 16580 20082 16646 20092
rect 16772 20082 16838 20092
rect 16964 20082 17030 20092
rect 17156 20082 17222 20092
rect 17348 20082 17414 20092
rect 17540 20082 17606 20092
rect 17732 20082 17798 20092
rect 17924 20082 17980 20092
rect 18408 20082 18474 20092
rect 18600 20082 18666 20092
rect 18792 20082 18858 20092
rect 18984 20082 19050 20092
rect 19176 20082 19242 20092
rect 19368 20082 19434 20092
rect 19560 20082 19626 20092
rect 19752 20082 19808 20092
rect 20236 20082 20302 20092
rect 20428 20082 20494 20092
rect 20620 20082 20686 20092
rect 20812 20082 20878 20092
rect 21004 20082 21070 20092
rect 21196 20082 21262 20092
rect 21388 20082 21454 20092
rect 21580 20082 21636 20092
rect 32 19744 98 19754
rect 224 19744 290 19754
rect 416 19744 482 19754
rect 608 19744 674 19754
rect 800 19744 866 19754
rect 992 19744 1058 19754
rect 1184 19744 1250 19754
rect 1376 19744 1442 19754
rect 1860 19744 1926 19754
rect 2052 19744 2118 19754
rect 2244 19744 2310 19754
rect 2436 19744 2502 19754
rect 2628 19744 2694 19754
rect 2820 19744 2886 19754
rect 3012 19744 3078 19754
rect 3204 19744 3270 19754
rect 3688 19744 3754 19754
rect 3880 19744 3946 19754
rect 4072 19744 4138 19754
rect 4264 19744 4330 19754
rect 4456 19744 4522 19754
rect 4648 19744 4714 19754
rect 4840 19744 4906 19754
rect 5032 19744 5098 19754
rect 5516 19744 5582 19754
rect 5708 19744 5774 19754
rect 5900 19744 5966 19754
rect 6092 19744 6158 19754
rect 6284 19744 6350 19754
rect 6476 19744 6542 19754
rect 6668 19744 6734 19754
rect 6860 19744 6926 19754
rect 7344 19744 7410 19754
rect 7536 19744 7602 19754
rect 7728 19744 7794 19754
rect 7920 19744 7986 19754
rect 8112 19744 8178 19754
rect 8304 19744 8370 19754
rect 8496 19744 8562 19754
rect 8688 19744 8754 19754
rect 9172 19744 9238 19754
rect 9364 19744 9430 19754
rect 9556 19744 9622 19754
rect 9748 19744 9814 19754
rect 9940 19744 10006 19754
rect 10132 19744 10198 19754
rect 10324 19744 10390 19754
rect 10516 19744 10582 19754
rect 11000 19744 11066 19754
rect 11192 19744 11258 19754
rect 11384 19744 11450 19754
rect 11576 19744 11642 19754
rect 11768 19744 11834 19754
rect 11960 19744 12026 19754
rect 12152 19744 12218 19754
rect 12344 19744 12410 19754
rect 12828 19744 12894 19754
rect 13020 19744 13086 19754
rect 13212 19744 13278 19754
rect 13404 19744 13470 19754
rect 13596 19744 13662 19754
rect 13788 19744 13854 19754
rect 13980 19744 14046 19754
rect 14172 19744 14238 19754
rect 14656 19744 14722 19754
rect 14848 19744 14914 19754
rect 15040 19744 15106 19754
rect 15232 19744 15298 19754
rect 15424 19744 15490 19754
rect 15616 19744 15682 19754
rect 15808 19744 15874 19754
rect 16000 19744 16066 19754
rect 16484 19744 16550 19754
rect 16676 19744 16742 19754
rect 16868 19744 16934 19754
rect 17060 19744 17126 19754
rect 17252 19744 17318 19754
rect 17444 19744 17510 19754
rect 17636 19744 17702 19754
rect 17828 19744 17894 19754
rect 18312 19744 18378 19754
rect 18504 19744 18570 19754
rect 18696 19744 18762 19754
rect 18888 19744 18954 19754
rect 19080 19744 19146 19754
rect 19272 19744 19338 19754
rect 19464 19744 19530 19754
rect 19656 19744 19722 19754
rect 20140 19744 20206 19754
rect 20332 19744 20398 19754
rect 20524 19744 20590 19754
rect 20716 19744 20782 19754
rect 20908 19744 20974 19754
rect 21100 19744 21166 19754
rect 21292 19744 21358 19754
rect 21484 19744 21550 19754
rect 0 19591 32 19744
rect 98 19591 224 19744
rect 290 19591 416 19744
rect 482 19591 608 19744
rect 674 19591 800 19744
rect 866 19591 992 19744
rect 1058 19591 1184 19744
rect 1250 19591 1376 19744
rect 1828 19591 1860 19744
rect 1926 19591 2052 19744
rect 2118 19591 2244 19744
rect 2310 19591 2436 19744
rect 2502 19591 2628 19744
rect 2694 19591 2820 19744
rect 2886 19591 3012 19744
rect 3078 19591 3204 19744
rect 3656 19591 3688 19744
rect 3754 19591 3880 19744
rect 3946 19591 4072 19744
rect 4138 19591 4264 19744
rect 4330 19591 4456 19744
rect 4522 19591 4648 19744
rect 4714 19591 4840 19744
rect 4906 19591 5032 19744
rect 5484 19591 5516 19744
rect 5582 19591 5708 19744
rect 5774 19591 5900 19744
rect 5966 19591 6092 19744
rect 6158 19591 6284 19744
rect 6350 19591 6476 19744
rect 6542 19591 6668 19744
rect 6734 19591 6860 19744
rect 7312 19591 7344 19744
rect 7410 19591 7536 19744
rect 7602 19591 7728 19744
rect 7794 19591 7920 19744
rect 7986 19591 8112 19744
rect 8178 19591 8304 19744
rect 8370 19591 8496 19744
rect 8562 19591 8688 19744
rect 9140 19591 9172 19744
rect 9238 19591 9364 19744
rect 9430 19591 9556 19744
rect 9622 19591 9748 19744
rect 9814 19591 9940 19744
rect 10006 19591 10132 19744
rect 10198 19591 10324 19744
rect 10390 19591 10516 19744
rect 10968 19591 11000 19744
rect 11066 19591 11192 19744
rect 11258 19591 11384 19744
rect 11450 19591 11576 19744
rect 11642 19591 11768 19744
rect 11834 19591 11960 19744
rect 12026 19591 12152 19744
rect 12218 19591 12344 19744
rect 12796 19591 12828 19744
rect 12894 19591 13020 19744
rect 13086 19591 13212 19744
rect 13278 19591 13404 19744
rect 13470 19591 13596 19744
rect 13662 19591 13788 19744
rect 13854 19591 13980 19744
rect 14046 19591 14172 19744
rect 14624 19591 14656 19744
rect 14722 19591 14848 19744
rect 14914 19591 15040 19744
rect 15106 19591 15232 19744
rect 15298 19591 15424 19744
rect 15490 19591 15616 19744
rect 15682 19591 15808 19744
rect 15874 19591 16000 19744
rect 16452 19591 16484 19744
rect 16550 19591 16676 19744
rect 16742 19591 16868 19744
rect 16934 19591 17060 19744
rect 17126 19591 17252 19744
rect 17318 19591 17444 19744
rect 17510 19591 17636 19744
rect 17702 19591 17828 19744
rect 18280 19591 18312 19744
rect 18378 19591 18504 19744
rect 18570 19591 18696 19744
rect 18762 19591 18888 19744
rect 18954 19591 19080 19744
rect 19146 19591 19272 19744
rect 19338 19591 19464 19744
rect 19530 19591 19656 19744
rect 20108 19591 20140 19744
rect 20206 19591 20332 19744
rect 20398 19591 20524 19744
rect 20590 19591 20716 19744
rect 20782 19591 20908 19744
rect 20974 19591 21100 19744
rect 21166 19591 21292 19744
rect 21358 19591 21484 19744
rect 32 19581 98 19591
rect 224 19581 290 19591
rect 416 19581 482 19591
rect 608 19581 674 19591
rect 800 19581 866 19591
rect 992 19581 1058 19591
rect 1184 19581 1250 19591
rect 1376 19581 1442 19591
rect 1860 19581 1926 19591
rect 2052 19581 2118 19591
rect 2244 19581 2310 19591
rect 2436 19581 2502 19591
rect 2628 19581 2694 19591
rect 2820 19581 2886 19591
rect 3012 19581 3078 19591
rect 3204 19581 3270 19591
rect 3688 19581 3754 19591
rect 3880 19581 3946 19591
rect 4072 19581 4138 19591
rect 4264 19581 4330 19591
rect 4456 19581 4522 19591
rect 4648 19581 4714 19591
rect 4840 19581 4906 19591
rect 5032 19581 5098 19591
rect 5516 19581 5582 19591
rect 5708 19581 5774 19591
rect 5900 19581 5966 19591
rect 6092 19581 6158 19591
rect 6284 19581 6350 19591
rect 6476 19581 6542 19591
rect 6668 19581 6734 19591
rect 6860 19581 6926 19591
rect 7344 19581 7410 19591
rect 7536 19581 7602 19591
rect 7728 19581 7794 19591
rect 7920 19581 7986 19591
rect 8112 19581 8178 19591
rect 8304 19581 8370 19591
rect 8496 19581 8562 19591
rect 8688 19581 8754 19591
rect 9172 19581 9238 19591
rect 9364 19581 9430 19591
rect 9556 19581 9622 19591
rect 9748 19581 9814 19591
rect 9940 19581 10006 19591
rect 10132 19581 10198 19591
rect 10324 19581 10390 19591
rect 10516 19581 10582 19591
rect 11000 19581 11066 19591
rect 11192 19581 11258 19591
rect 11384 19581 11450 19591
rect 11576 19581 11642 19591
rect 11768 19581 11834 19591
rect 11960 19581 12026 19591
rect 12152 19581 12218 19591
rect 12344 19581 12410 19591
rect 12828 19581 12894 19591
rect 13020 19581 13086 19591
rect 13212 19581 13278 19591
rect 13404 19581 13470 19591
rect 13596 19581 13662 19591
rect 13788 19581 13854 19591
rect 13980 19581 14046 19591
rect 14172 19581 14238 19591
rect 14656 19581 14722 19591
rect 14848 19581 14914 19591
rect 15040 19581 15106 19591
rect 15232 19581 15298 19591
rect 15424 19581 15490 19591
rect 15616 19581 15682 19591
rect 15808 19581 15874 19591
rect 16000 19581 16066 19591
rect 16484 19581 16550 19591
rect 16676 19581 16742 19591
rect 16868 19581 16934 19591
rect 17060 19581 17126 19591
rect 17252 19581 17318 19591
rect 17444 19581 17510 19591
rect 17636 19581 17702 19591
rect 17828 19581 17894 19591
rect 18312 19581 18378 19591
rect 18504 19581 18570 19591
rect 18696 19581 18762 19591
rect 18888 19581 18954 19591
rect 19080 19581 19146 19591
rect 19272 19581 19338 19591
rect 19464 19581 19530 19591
rect 19656 19581 19722 19591
rect 20140 19581 20206 19591
rect 20332 19581 20398 19591
rect 20524 19581 20590 19591
rect 20716 19581 20782 19591
rect 20908 19581 20974 19591
rect 21100 19581 21166 19591
rect 21292 19581 21358 19591
rect 21484 19581 21550 19591
rect 128 19531 194 19541
rect 320 19531 386 19541
rect 512 19531 578 19541
rect 704 19531 770 19541
rect 896 19531 962 19541
rect 1088 19531 1154 19541
rect 1280 19531 1346 19541
rect 1472 19531 1528 19541
rect 1956 19531 2022 19541
rect 2148 19531 2214 19541
rect 2340 19531 2406 19541
rect 2532 19531 2598 19541
rect 2724 19531 2790 19541
rect 2916 19531 2982 19541
rect 3108 19531 3174 19541
rect 3300 19531 3356 19541
rect 3784 19531 3850 19541
rect 3976 19531 4042 19541
rect 4168 19531 4234 19541
rect 4360 19531 4426 19541
rect 4552 19531 4618 19541
rect 4744 19531 4810 19541
rect 4936 19531 5002 19541
rect 5128 19531 5184 19541
rect 5612 19531 5678 19541
rect 5804 19531 5870 19541
rect 5996 19531 6062 19541
rect 6188 19531 6254 19541
rect 6380 19531 6446 19541
rect 6572 19531 6638 19541
rect 6764 19531 6830 19541
rect 6956 19531 7012 19541
rect 7440 19531 7506 19541
rect 7632 19531 7698 19541
rect 7824 19531 7890 19541
rect 8016 19531 8082 19541
rect 8208 19531 8274 19541
rect 8400 19531 8466 19541
rect 8592 19531 8658 19541
rect 8784 19531 8840 19541
rect 9268 19531 9334 19541
rect 9460 19531 9526 19541
rect 9652 19531 9718 19541
rect 9844 19531 9910 19541
rect 10036 19531 10102 19541
rect 10228 19531 10294 19541
rect 10420 19531 10486 19541
rect 10612 19531 10668 19541
rect 11096 19531 11162 19541
rect 11288 19531 11354 19541
rect 11480 19531 11546 19541
rect 11672 19531 11738 19541
rect 11864 19531 11930 19541
rect 12056 19531 12122 19541
rect 12248 19531 12314 19541
rect 12440 19531 12496 19541
rect 12924 19531 12990 19541
rect 13116 19531 13182 19541
rect 13308 19531 13374 19541
rect 13500 19531 13566 19541
rect 13692 19531 13758 19541
rect 13884 19531 13950 19541
rect 14076 19531 14142 19541
rect 14268 19531 14324 19541
rect 14752 19531 14818 19541
rect 14944 19531 15010 19541
rect 15136 19531 15202 19541
rect 15328 19531 15394 19541
rect 15520 19531 15586 19541
rect 15712 19531 15778 19541
rect 15904 19531 15970 19541
rect 16096 19531 16152 19541
rect 16580 19531 16646 19541
rect 16772 19531 16838 19541
rect 16964 19531 17030 19541
rect 17156 19531 17222 19541
rect 17348 19531 17414 19541
rect 17540 19531 17606 19541
rect 17732 19531 17798 19541
rect 17924 19531 17980 19541
rect 18408 19531 18474 19541
rect 18600 19531 18666 19541
rect 18792 19531 18858 19541
rect 18984 19531 19050 19541
rect 19176 19531 19242 19541
rect 19368 19531 19434 19541
rect 19560 19531 19626 19541
rect 19752 19531 19808 19541
rect 20236 19531 20302 19541
rect 20428 19531 20494 19541
rect 20620 19531 20686 19541
rect 20812 19531 20878 19541
rect 21004 19531 21070 19541
rect 21196 19531 21262 19541
rect 21388 19531 21454 19541
rect 21580 19531 21636 19541
rect 0 19378 128 19531
rect 194 19378 320 19531
rect 386 19378 512 19531
rect 578 19378 704 19531
rect 770 19378 896 19531
rect 962 19378 1088 19531
rect 1154 19378 1280 19531
rect 1346 19378 1472 19531
rect 1528 19378 1708 19531
rect 1828 19378 1956 19531
rect 2022 19378 2148 19531
rect 2214 19378 2340 19531
rect 2406 19378 2532 19531
rect 2598 19378 2724 19531
rect 2790 19378 2916 19531
rect 2982 19378 3108 19531
rect 3174 19378 3300 19531
rect 3356 19378 3536 19531
rect 3656 19378 3784 19531
rect 3850 19378 3976 19531
rect 4042 19378 4168 19531
rect 4234 19378 4360 19531
rect 4426 19378 4552 19531
rect 4618 19378 4744 19531
rect 4810 19378 4936 19531
rect 5002 19378 5128 19531
rect 5184 19378 5364 19531
rect 5484 19378 5612 19531
rect 5678 19378 5804 19531
rect 5870 19378 5996 19531
rect 6062 19378 6188 19531
rect 6254 19378 6380 19531
rect 6446 19378 6572 19531
rect 6638 19378 6764 19531
rect 6830 19378 6956 19531
rect 7012 19378 7192 19531
rect 7312 19378 7440 19531
rect 7506 19378 7632 19531
rect 7698 19378 7824 19531
rect 7890 19378 8016 19531
rect 8082 19378 8208 19531
rect 8274 19378 8400 19531
rect 8466 19378 8592 19531
rect 8658 19378 8784 19531
rect 8840 19378 9020 19531
rect 9140 19378 9268 19531
rect 9334 19378 9460 19531
rect 9526 19378 9652 19531
rect 9718 19378 9844 19531
rect 9910 19378 10036 19531
rect 10102 19378 10228 19531
rect 10294 19378 10420 19531
rect 10486 19378 10612 19531
rect 10668 19378 10848 19531
rect 10968 19378 11096 19531
rect 11162 19378 11288 19531
rect 11354 19378 11480 19531
rect 11546 19378 11672 19531
rect 11738 19378 11864 19531
rect 11930 19378 12056 19531
rect 12122 19378 12248 19531
rect 12314 19378 12440 19531
rect 12496 19378 12676 19531
rect 12796 19378 12924 19531
rect 12990 19378 13116 19531
rect 13182 19378 13308 19531
rect 13374 19378 13500 19531
rect 13566 19378 13692 19531
rect 13758 19378 13884 19531
rect 13950 19378 14076 19531
rect 14142 19378 14268 19531
rect 14324 19378 14504 19531
rect 14624 19378 14752 19531
rect 14818 19378 14944 19531
rect 15010 19378 15136 19531
rect 15202 19378 15328 19531
rect 15394 19378 15520 19531
rect 15586 19378 15712 19531
rect 15778 19378 15904 19531
rect 15970 19378 16096 19531
rect 16152 19378 16332 19531
rect 16452 19378 16580 19531
rect 16646 19378 16772 19531
rect 16838 19378 16964 19531
rect 17030 19378 17156 19531
rect 17222 19378 17348 19531
rect 17414 19378 17540 19531
rect 17606 19378 17732 19531
rect 17798 19378 17924 19531
rect 17980 19378 18160 19531
rect 18280 19378 18408 19531
rect 18474 19378 18600 19531
rect 18666 19378 18792 19531
rect 18858 19378 18984 19531
rect 19050 19378 19176 19531
rect 19242 19378 19368 19531
rect 19434 19378 19560 19531
rect 19626 19378 19752 19531
rect 19808 19378 19988 19531
rect 20108 19378 20236 19531
rect 20302 19378 20428 19531
rect 20494 19378 20620 19531
rect 20686 19378 20812 19531
rect 20878 19378 21004 19531
rect 21070 19378 21196 19531
rect 21262 19378 21388 19531
rect 21454 19378 21580 19531
rect 21636 19378 21816 19531
rect 128 19368 194 19378
rect 320 19368 386 19378
rect 512 19368 578 19378
rect 704 19368 770 19378
rect 896 19368 962 19378
rect 1088 19368 1154 19378
rect 1280 19368 1346 19378
rect 1472 19368 1528 19378
rect 1956 19368 2022 19378
rect 2148 19368 2214 19378
rect 2340 19368 2406 19378
rect 2532 19368 2598 19378
rect 2724 19368 2790 19378
rect 2916 19368 2982 19378
rect 3108 19368 3174 19378
rect 3300 19368 3356 19378
rect 3784 19368 3850 19378
rect 3976 19368 4042 19378
rect 4168 19368 4234 19378
rect 4360 19368 4426 19378
rect 4552 19368 4618 19378
rect 4744 19368 4810 19378
rect 4936 19368 5002 19378
rect 5128 19368 5184 19378
rect 5612 19368 5678 19378
rect 5804 19368 5870 19378
rect 5996 19368 6062 19378
rect 6188 19368 6254 19378
rect 6380 19368 6446 19378
rect 6572 19368 6638 19378
rect 6764 19368 6830 19378
rect 6956 19368 7012 19378
rect 7440 19368 7506 19378
rect 7632 19368 7698 19378
rect 7824 19368 7890 19378
rect 8016 19368 8082 19378
rect 8208 19368 8274 19378
rect 8400 19368 8466 19378
rect 8592 19368 8658 19378
rect 8784 19368 8840 19378
rect 9268 19368 9334 19378
rect 9460 19368 9526 19378
rect 9652 19368 9718 19378
rect 9844 19368 9910 19378
rect 10036 19368 10102 19378
rect 10228 19368 10294 19378
rect 10420 19368 10486 19378
rect 10612 19368 10668 19378
rect 11096 19368 11162 19378
rect 11288 19368 11354 19378
rect 11480 19368 11546 19378
rect 11672 19368 11738 19378
rect 11864 19368 11930 19378
rect 12056 19368 12122 19378
rect 12248 19368 12314 19378
rect 12440 19368 12496 19378
rect 12924 19368 12990 19378
rect 13116 19368 13182 19378
rect 13308 19368 13374 19378
rect 13500 19368 13566 19378
rect 13692 19368 13758 19378
rect 13884 19368 13950 19378
rect 14076 19368 14142 19378
rect 14268 19368 14324 19378
rect 14752 19368 14818 19378
rect 14944 19368 15010 19378
rect 15136 19368 15202 19378
rect 15328 19368 15394 19378
rect 15520 19368 15586 19378
rect 15712 19368 15778 19378
rect 15904 19368 15970 19378
rect 16096 19368 16152 19378
rect 16580 19368 16646 19378
rect 16772 19368 16838 19378
rect 16964 19368 17030 19378
rect 17156 19368 17222 19378
rect 17348 19368 17414 19378
rect 17540 19368 17606 19378
rect 17732 19368 17798 19378
rect 17924 19368 17980 19378
rect 18408 19368 18474 19378
rect 18600 19368 18666 19378
rect 18792 19368 18858 19378
rect 18984 19368 19050 19378
rect 19176 19368 19242 19378
rect 19368 19368 19434 19378
rect 19560 19368 19626 19378
rect 19752 19368 19808 19378
rect 20236 19368 20302 19378
rect 20428 19368 20494 19378
rect 20620 19368 20686 19378
rect 20812 19368 20878 19378
rect 21004 19368 21070 19378
rect 21196 19368 21262 19378
rect 21388 19368 21454 19378
rect 21580 19368 21636 19378
rect 32 19030 98 19040
rect 224 19030 290 19040
rect 416 19030 482 19040
rect 608 19030 674 19040
rect 800 19030 866 19040
rect 992 19030 1058 19040
rect 1184 19030 1250 19040
rect 1376 19030 1442 19040
rect 1860 19030 1926 19040
rect 2052 19030 2118 19040
rect 2244 19030 2310 19040
rect 2436 19030 2502 19040
rect 2628 19030 2694 19040
rect 2820 19030 2886 19040
rect 3012 19030 3078 19040
rect 3204 19030 3270 19040
rect 3688 19030 3754 19040
rect 3880 19030 3946 19040
rect 4072 19030 4138 19040
rect 4264 19030 4330 19040
rect 4456 19030 4522 19040
rect 4648 19030 4714 19040
rect 4840 19030 4906 19040
rect 5032 19030 5098 19040
rect 5516 19030 5582 19040
rect 5708 19030 5774 19040
rect 5900 19030 5966 19040
rect 6092 19030 6158 19040
rect 6284 19030 6350 19040
rect 6476 19030 6542 19040
rect 6668 19030 6734 19040
rect 6860 19030 6926 19040
rect 7344 19030 7410 19040
rect 7536 19030 7602 19040
rect 7728 19030 7794 19040
rect 7920 19030 7986 19040
rect 8112 19030 8178 19040
rect 8304 19030 8370 19040
rect 8496 19030 8562 19040
rect 8688 19030 8754 19040
rect 9172 19030 9238 19040
rect 9364 19030 9430 19040
rect 9556 19030 9622 19040
rect 9748 19030 9814 19040
rect 9940 19030 10006 19040
rect 10132 19030 10198 19040
rect 10324 19030 10390 19040
rect 10516 19030 10582 19040
rect 11000 19030 11066 19040
rect 11192 19030 11258 19040
rect 11384 19030 11450 19040
rect 11576 19030 11642 19040
rect 11768 19030 11834 19040
rect 11960 19030 12026 19040
rect 12152 19030 12218 19040
rect 12344 19030 12410 19040
rect 12828 19030 12894 19040
rect 13020 19030 13086 19040
rect 13212 19030 13278 19040
rect 13404 19030 13470 19040
rect 13596 19030 13662 19040
rect 13788 19030 13854 19040
rect 13980 19030 14046 19040
rect 14172 19030 14238 19040
rect 14656 19030 14722 19040
rect 14848 19030 14914 19040
rect 15040 19030 15106 19040
rect 15232 19030 15298 19040
rect 15424 19030 15490 19040
rect 15616 19030 15682 19040
rect 15808 19030 15874 19040
rect 16000 19030 16066 19040
rect 16484 19030 16550 19040
rect 16676 19030 16742 19040
rect 16868 19030 16934 19040
rect 17060 19030 17126 19040
rect 17252 19030 17318 19040
rect 17444 19030 17510 19040
rect 17636 19030 17702 19040
rect 17828 19030 17894 19040
rect 18312 19030 18378 19040
rect 18504 19030 18570 19040
rect 18696 19030 18762 19040
rect 18888 19030 18954 19040
rect 19080 19030 19146 19040
rect 19272 19030 19338 19040
rect 19464 19030 19530 19040
rect 19656 19030 19722 19040
rect 20140 19030 20206 19040
rect 20332 19030 20398 19040
rect 20524 19030 20590 19040
rect 20716 19030 20782 19040
rect 20908 19030 20974 19040
rect 21100 19030 21166 19040
rect 21292 19030 21358 19040
rect 21484 19030 21550 19040
rect 0 18877 32 19030
rect 98 18877 224 19030
rect 290 18877 416 19030
rect 482 18877 608 19030
rect 674 18877 800 19030
rect 866 18877 992 19030
rect 1058 18877 1184 19030
rect 1250 18877 1376 19030
rect 1828 18877 1860 19030
rect 1926 18877 2052 19030
rect 2118 18877 2244 19030
rect 2310 18877 2436 19030
rect 2502 18877 2628 19030
rect 2694 18877 2820 19030
rect 2886 18877 3012 19030
rect 3078 18877 3204 19030
rect 3656 18877 3688 19030
rect 3754 18877 3880 19030
rect 3946 18877 4072 19030
rect 4138 18877 4264 19030
rect 4330 18877 4456 19030
rect 4522 18877 4648 19030
rect 4714 18877 4840 19030
rect 4906 18877 5032 19030
rect 5484 18877 5516 19030
rect 5582 18877 5708 19030
rect 5774 18877 5900 19030
rect 5966 18877 6092 19030
rect 6158 18877 6284 19030
rect 6350 18877 6476 19030
rect 6542 18877 6668 19030
rect 6734 18877 6860 19030
rect 7312 18877 7344 19030
rect 7410 18877 7536 19030
rect 7602 18877 7728 19030
rect 7794 18877 7920 19030
rect 7986 18877 8112 19030
rect 8178 18877 8304 19030
rect 8370 18877 8496 19030
rect 8562 18877 8688 19030
rect 9140 18877 9172 19030
rect 9238 18877 9364 19030
rect 9430 18877 9556 19030
rect 9622 18877 9748 19030
rect 9814 18877 9940 19030
rect 10006 18877 10132 19030
rect 10198 18877 10324 19030
rect 10390 18877 10516 19030
rect 10968 18877 11000 19030
rect 11066 18877 11192 19030
rect 11258 18877 11384 19030
rect 11450 18877 11576 19030
rect 11642 18877 11768 19030
rect 11834 18877 11960 19030
rect 12026 18877 12152 19030
rect 12218 18877 12344 19030
rect 12796 18877 12828 19030
rect 12894 18877 13020 19030
rect 13086 18877 13212 19030
rect 13278 18877 13404 19030
rect 13470 18877 13596 19030
rect 13662 18877 13788 19030
rect 13854 18877 13980 19030
rect 14046 18877 14172 19030
rect 14624 18877 14656 19030
rect 14722 18877 14848 19030
rect 14914 18877 15040 19030
rect 15106 18877 15232 19030
rect 15298 18877 15424 19030
rect 15490 18877 15616 19030
rect 15682 18877 15808 19030
rect 15874 18877 16000 19030
rect 16452 18877 16484 19030
rect 16550 18877 16676 19030
rect 16742 18877 16868 19030
rect 16934 18877 17060 19030
rect 17126 18877 17252 19030
rect 17318 18877 17444 19030
rect 17510 18877 17636 19030
rect 17702 18877 17828 19030
rect 18280 18877 18312 19030
rect 18378 18877 18504 19030
rect 18570 18877 18696 19030
rect 18762 18877 18888 19030
rect 18954 18877 19080 19030
rect 19146 18877 19272 19030
rect 19338 18877 19464 19030
rect 19530 18877 19656 19030
rect 20108 18877 20140 19030
rect 20206 18877 20332 19030
rect 20398 18877 20524 19030
rect 20590 18877 20716 19030
rect 20782 18877 20908 19030
rect 20974 18877 21100 19030
rect 21166 18877 21292 19030
rect 21358 18877 21484 19030
rect 32 18867 98 18877
rect 224 18867 290 18877
rect 416 18867 482 18877
rect 608 18867 674 18877
rect 800 18867 866 18877
rect 992 18867 1058 18877
rect 1184 18867 1250 18877
rect 1376 18867 1442 18877
rect 1860 18867 1926 18877
rect 2052 18867 2118 18877
rect 2244 18867 2310 18877
rect 2436 18867 2502 18877
rect 2628 18867 2694 18877
rect 2820 18867 2886 18877
rect 3012 18867 3078 18877
rect 3204 18867 3270 18877
rect 3688 18867 3754 18877
rect 3880 18867 3946 18877
rect 4072 18867 4138 18877
rect 4264 18867 4330 18877
rect 4456 18867 4522 18877
rect 4648 18867 4714 18877
rect 4840 18867 4906 18877
rect 5032 18867 5098 18877
rect 5516 18867 5582 18877
rect 5708 18867 5774 18877
rect 5900 18867 5966 18877
rect 6092 18867 6158 18877
rect 6284 18867 6350 18877
rect 6476 18867 6542 18877
rect 6668 18867 6734 18877
rect 6860 18867 6926 18877
rect 7344 18867 7410 18877
rect 7536 18867 7602 18877
rect 7728 18867 7794 18877
rect 7920 18867 7986 18877
rect 8112 18867 8178 18877
rect 8304 18867 8370 18877
rect 8496 18867 8562 18877
rect 8688 18867 8754 18877
rect 9172 18867 9238 18877
rect 9364 18867 9430 18877
rect 9556 18867 9622 18877
rect 9748 18867 9814 18877
rect 9940 18867 10006 18877
rect 10132 18867 10198 18877
rect 10324 18867 10390 18877
rect 10516 18867 10582 18877
rect 11000 18867 11066 18877
rect 11192 18867 11258 18877
rect 11384 18867 11450 18877
rect 11576 18867 11642 18877
rect 11768 18867 11834 18877
rect 11960 18867 12026 18877
rect 12152 18867 12218 18877
rect 12344 18867 12410 18877
rect 12828 18867 12894 18877
rect 13020 18867 13086 18877
rect 13212 18867 13278 18877
rect 13404 18867 13470 18877
rect 13596 18867 13662 18877
rect 13788 18867 13854 18877
rect 13980 18867 14046 18877
rect 14172 18867 14238 18877
rect 14656 18867 14722 18877
rect 14848 18867 14914 18877
rect 15040 18867 15106 18877
rect 15232 18867 15298 18877
rect 15424 18867 15490 18877
rect 15616 18867 15682 18877
rect 15808 18867 15874 18877
rect 16000 18867 16066 18877
rect 16484 18867 16550 18877
rect 16676 18867 16742 18877
rect 16868 18867 16934 18877
rect 17060 18867 17126 18877
rect 17252 18867 17318 18877
rect 17444 18867 17510 18877
rect 17636 18867 17702 18877
rect 17828 18867 17894 18877
rect 18312 18867 18378 18877
rect 18504 18867 18570 18877
rect 18696 18867 18762 18877
rect 18888 18867 18954 18877
rect 19080 18867 19146 18877
rect 19272 18867 19338 18877
rect 19464 18867 19530 18877
rect 19656 18867 19722 18877
rect 20140 18867 20206 18877
rect 20332 18867 20398 18877
rect 20524 18867 20590 18877
rect 20716 18867 20782 18877
rect 20908 18867 20974 18877
rect 21100 18867 21166 18877
rect 21292 18867 21358 18877
rect 21484 18867 21550 18877
rect 128 18817 194 18827
rect 320 18817 386 18827
rect 512 18817 578 18827
rect 704 18817 770 18827
rect 896 18817 962 18827
rect 1088 18817 1154 18827
rect 1280 18817 1346 18827
rect 1472 18817 1528 18827
rect 1956 18817 2022 18827
rect 2148 18817 2214 18827
rect 2340 18817 2406 18827
rect 2532 18817 2598 18827
rect 2724 18817 2790 18827
rect 2916 18817 2982 18827
rect 3108 18817 3174 18827
rect 3300 18817 3356 18827
rect 3784 18817 3850 18827
rect 3976 18817 4042 18827
rect 4168 18817 4234 18827
rect 4360 18817 4426 18827
rect 4552 18817 4618 18827
rect 4744 18817 4810 18827
rect 4936 18817 5002 18827
rect 5128 18817 5184 18827
rect 5612 18817 5678 18827
rect 5804 18817 5870 18827
rect 5996 18817 6062 18827
rect 6188 18817 6254 18827
rect 6380 18817 6446 18827
rect 6572 18817 6638 18827
rect 6764 18817 6830 18827
rect 6956 18817 7012 18827
rect 7440 18817 7506 18827
rect 7632 18817 7698 18827
rect 7824 18817 7890 18827
rect 8016 18817 8082 18827
rect 8208 18817 8274 18827
rect 8400 18817 8466 18827
rect 8592 18817 8658 18827
rect 8784 18817 8840 18827
rect 9268 18817 9334 18827
rect 9460 18817 9526 18827
rect 9652 18817 9718 18827
rect 9844 18817 9910 18827
rect 10036 18817 10102 18827
rect 10228 18817 10294 18827
rect 10420 18817 10486 18827
rect 10612 18817 10668 18827
rect 11096 18817 11162 18827
rect 11288 18817 11354 18827
rect 11480 18817 11546 18827
rect 11672 18817 11738 18827
rect 11864 18817 11930 18827
rect 12056 18817 12122 18827
rect 12248 18817 12314 18827
rect 12440 18817 12496 18827
rect 12924 18817 12990 18827
rect 13116 18817 13182 18827
rect 13308 18817 13374 18827
rect 13500 18817 13566 18827
rect 13692 18817 13758 18827
rect 13884 18817 13950 18827
rect 14076 18817 14142 18827
rect 14268 18817 14324 18827
rect 14752 18817 14818 18827
rect 14944 18817 15010 18827
rect 15136 18817 15202 18827
rect 15328 18817 15394 18827
rect 15520 18817 15586 18827
rect 15712 18817 15778 18827
rect 15904 18817 15970 18827
rect 16096 18817 16152 18827
rect 16580 18817 16646 18827
rect 16772 18817 16838 18827
rect 16964 18817 17030 18827
rect 17156 18817 17222 18827
rect 17348 18817 17414 18827
rect 17540 18817 17606 18827
rect 17732 18817 17798 18827
rect 17924 18817 17980 18827
rect 18408 18817 18474 18827
rect 18600 18817 18666 18827
rect 18792 18817 18858 18827
rect 18984 18817 19050 18827
rect 19176 18817 19242 18827
rect 19368 18817 19434 18827
rect 19560 18817 19626 18827
rect 19752 18817 19808 18827
rect 20236 18817 20302 18827
rect 20428 18817 20494 18827
rect 20620 18817 20686 18827
rect 20812 18817 20878 18827
rect 21004 18817 21070 18827
rect 21196 18817 21262 18827
rect 21388 18817 21454 18827
rect 21580 18817 21636 18827
rect 0 18664 128 18817
rect 194 18664 320 18817
rect 386 18664 512 18817
rect 578 18664 704 18817
rect 770 18664 896 18817
rect 962 18664 1088 18817
rect 1154 18664 1280 18817
rect 1346 18664 1472 18817
rect 1528 18664 1708 18817
rect 1828 18664 1956 18817
rect 2022 18664 2148 18817
rect 2214 18664 2340 18817
rect 2406 18664 2532 18817
rect 2598 18664 2724 18817
rect 2790 18664 2916 18817
rect 2982 18664 3108 18817
rect 3174 18664 3300 18817
rect 3356 18664 3536 18817
rect 3656 18664 3784 18817
rect 3850 18664 3976 18817
rect 4042 18664 4168 18817
rect 4234 18664 4360 18817
rect 4426 18664 4552 18817
rect 4618 18664 4744 18817
rect 4810 18664 4936 18817
rect 5002 18664 5128 18817
rect 5184 18664 5364 18817
rect 5484 18664 5612 18817
rect 5678 18664 5804 18817
rect 5870 18664 5996 18817
rect 6062 18664 6188 18817
rect 6254 18664 6380 18817
rect 6446 18664 6572 18817
rect 6638 18664 6764 18817
rect 6830 18664 6956 18817
rect 7012 18664 7192 18817
rect 7312 18664 7440 18817
rect 7506 18664 7632 18817
rect 7698 18664 7824 18817
rect 7890 18664 8016 18817
rect 8082 18664 8208 18817
rect 8274 18664 8400 18817
rect 8466 18664 8592 18817
rect 8658 18664 8784 18817
rect 8840 18664 9020 18817
rect 9140 18664 9268 18817
rect 9334 18664 9460 18817
rect 9526 18664 9652 18817
rect 9718 18664 9844 18817
rect 9910 18664 10036 18817
rect 10102 18664 10228 18817
rect 10294 18664 10420 18817
rect 10486 18664 10612 18817
rect 10668 18664 10848 18817
rect 10968 18664 11096 18817
rect 11162 18664 11288 18817
rect 11354 18664 11480 18817
rect 11546 18664 11672 18817
rect 11738 18664 11864 18817
rect 11930 18664 12056 18817
rect 12122 18664 12248 18817
rect 12314 18664 12440 18817
rect 12496 18664 12676 18817
rect 12796 18664 12924 18817
rect 12990 18664 13116 18817
rect 13182 18664 13308 18817
rect 13374 18664 13500 18817
rect 13566 18664 13692 18817
rect 13758 18664 13884 18817
rect 13950 18664 14076 18817
rect 14142 18664 14268 18817
rect 14324 18664 14504 18817
rect 14624 18664 14752 18817
rect 14818 18664 14944 18817
rect 15010 18664 15136 18817
rect 15202 18664 15328 18817
rect 15394 18664 15520 18817
rect 15586 18664 15712 18817
rect 15778 18664 15904 18817
rect 15970 18664 16096 18817
rect 16152 18664 16332 18817
rect 16452 18664 16580 18817
rect 16646 18664 16772 18817
rect 16838 18664 16964 18817
rect 17030 18664 17156 18817
rect 17222 18664 17348 18817
rect 17414 18664 17540 18817
rect 17606 18664 17732 18817
rect 17798 18664 17924 18817
rect 17980 18664 18160 18817
rect 18280 18664 18408 18817
rect 18474 18664 18600 18817
rect 18666 18664 18792 18817
rect 18858 18664 18984 18817
rect 19050 18664 19176 18817
rect 19242 18664 19368 18817
rect 19434 18664 19560 18817
rect 19626 18664 19752 18817
rect 19808 18664 19988 18817
rect 20108 18664 20236 18817
rect 20302 18664 20428 18817
rect 20494 18664 20620 18817
rect 20686 18664 20812 18817
rect 20878 18664 21004 18817
rect 21070 18664 21196 18817
rect 21262 18664 21388 18817
rect 21454 18664 21580 18817
rect 21636 18664 21816 18817
rect 128 18654 194 18664
rect 320 18654 386 18664
rect 512 18654 578 18664
rect 704 18654 770 18664
rect 896 18654 962 18664
rect 1088 18654 1154 18664
rect 1280 18654 1346 18664
rect 1472 18654 1528 18664
rect 1956 18654 2022 18664
rect 2148 18654 2214 18664
rect 2340 18654 2406 18664
rect 2532 18654 2598 18664
rect 2724 18654 2790 18664
rect 2916 18654 2982 18664
rect 3108 18654 3174 18664
rect 3300 18654 3356 18664
rect 3784 18654 3850 18664
rect 3976 18654 4042 18664
rect 4168 18654 4234 18664
rect 4360 18654 4426 18664
rect 4552 18654 4618 18664
rect 4744 18654 4810 18664
rect 4936 18654 5002 18664
rect 5128 18654 5184 18664
rect 5612 18654 5678 18664
rect 5804 18654 5870 18664
rect 5996 18654 6062 18664
rect 6188 18654 6254 18664
rect 6380 18654 6446 18664
rect 6572 18654 6638 18664
rect 6764 18654 6830 18664
rect 6956 18654 7012 18664
rect 7440 18654 7506 18664
rect 7632 18654 7698 18664
rect 7824 18654 7890 18664
rect 8016 18654 8082 18664
rect 8208 18654 8274 18664
rect 8400 18654 8466 18664
rect 8592 18654 8658 18664
rect 8784 18654 8840 18664
rect 9268 18654 9334 18664
rect 9460 18654 9526 18664
rect 9652 18654 9718 18664
rect 9844 18654 9910 18664
rect 10036 18654 10102 18664
rect 10228 18654 10294 18664
rect 10420 18654 10486 18664
rect 10612 18654 10668 18664
rect 11096 18654 11162 18664
rect 11288 18654 11354 18664
rect 11480 18654 11546 18664
rect 11672 18654 11738 18664
rect 11864 18654 11930 18664
rect 12056 18654 12122 18664
rect 12248 18654 12314 18664
rect 12440 18654 12496 18664
rect 12924 18654 12990 18664
rect 13116 18654 13182 18664
rect 13308 18654 13374 18664
rect 13500 18654 13566 18664
rect 13692 18654 13758 18664
rect 13884 18654 13950 18664
rect 14076 18654 14142 18664
rect 14268 18654 14324 18664
rect 14752 18654 14818 18664
rect 14944 18654 15010 18664
rect 15136 18654 15202 18664
rect 15328 18654 15394 18664
rect 15520 18654 15586 18664
rect 15712 18654 15778 18664
rect 15904 18654 15970 18664
rect 16096 18654 16152 18664
rect 16580 18654 16646 18664
rect 16772 18654 16838 18664
rect 16964 18654 17030 18664
rect 17156 18654 17222 18664
rect 17348 18654 17414 18664
rect 17540 18654 17606 18664
rect 17732 18654 17798 18664
rect 17924 18654 17980 18664
rect 18408 18654 18474 18664
rect 18600 18654 18666 18664
rect 18792 18654 18858 18664
rect 18984 18654 19050 18664
rect 19176 18654 19242 18664
rect 19368 18654 19434 18664
rect 19560 18654 19626 18664
rect 19752 18654 19808 18664
rect 20236 18654 20302 18664
rect 20428 18654 20494 18664
rect 20620 18654 20686 18664
rect 20812 18654 20878 18664
rect 21004 18654 21070 18664
rect 21196 18654 21262 18664
rect 21388 18654 21454 18664
rect 21580 18654 21636 18664
rect 32 18316 98 18326
rect 224 18316 290 18326
rect 416 18316 482 18326
rect 608 18316 674 18326
rect 800 18316 866 18326
rect 992 18316 1058 18326
rect 1184 18316 1250 18326
rect 1376 18316 1442 18326
rect 1860 18316 1926 18326
rect 2052 18316 2118 18326
rect 2244 18316 2310 18326
rect 2436 18316 2502 18326
rect 2628 18316 2694 18326
rect 2820 18316 2886 18326
rect 3012 18316 3078 18326
rect 3204 18316 3270 18326
rect 3688 18316 3754 18326
rect 3880 18316 3946 18326
rect 4072 18316 4138 18326
rect 4264 18316 4330 18326
rect 4456 18316 4522 18326
rect 4648 18316 4714 18326
rect 4840 18316 4906 18326
rect 5032 18316 5098 18326
rect 5516 18316 5582 18326
rect 5708 18316 5774 18326
rect 5900 18316 5966 18326
rect 6092 18316 6158 18326
rect 6284 18316 6350 18326
rect 6476 18316 6542 18326
rect 6668 18316 6734 18326
rect 6860 18316 6926 18326
rect 7344 18316 7410 18326
rect 7536 18316 7602 18326
rect 7728 18316 7794 18326
rect 7920 18316 7986 18326
rect 8112 18316 8178 18326
rect 8304 18316 8370 18326
rect 8496 18316 8562 18326
rect 8688 18316 8754 18326
rect 9172 18316 9238 18326
rect 9364 18316 9430 18326
rect 9556 18316 9622 18326
rect 9748 18316 9814 18326
rect 9940 18316 10006 18326
rect 10132 18316 10198 18326
rect 10324 18316 10390 18326
rect 10516 18316 10582 18326
rect 11000 18316 11066 18326
rect 11192 18316 11258 18326
rect 11384 18316 11450 18326
rect 11576 18316 11642 18326
rect 11768 18316 11834 18326
rect 11960 18316 12026 18326
rect 12152 18316 12218 18326
rect 12344 18316 12410 18326
rect 12828 18316 12894 18326
rect 13020 18316 13086 18326
rect 13212 18316 13278 18326
rect 13404 18316 13470 18326
rect 13596 18316 13662 18326
rect 13788 18316 13854 18326
rect 13980 18316 14046 18326
rect 14172 18316 14238 18326
rect 14656 18316 14722 18326
rect 14848 18316 14914 18326
rect 15040 18316 15106 18326
rect 15232 18316 15298 18326
rect 15424 18316 15490 18326
rect 15616 18316 15682 18326
rect 15808 18316 15874 18326
rect 16000 18316 16066 18326
rect 16484 18316 16550 18326
rect 16676 18316 16742 18326
rect 16868 18316 16934 18326
rect 17060 18316 17126 18326
rect 17252 18316 17318 18326
rect 17444 18316 17510 18326
rect 17636 18316 17702 18326
rect 17828 18316 17894 18326
rect 18312 18316 18378 18326
rect 18504 18316 18570 18326
rect 18696 18316 18762 18326
rect 18888 18316 18954 18326
rect 19080 18316 19146 18326
rect 19272 18316 19338 18326
rect 19464 18316 19530 18326
rect 19656 18316 19722 18326
rect 20140 18316 20206 18326
rect 20332 18316 20398 18326
rect 20524 18316 20590 18326
rect 20716 18316 20782 18326
rect 20908 18316 20974 18326
rect 21100 18316 21166 18326
rect 21292 18316 21358 18326
rect 21484 18316 21550 18326
rect 0 18163 32 18316
rect 98 18163 224 18316
rect 290 18163 416 18316
rect 482 18163 608 18316
rect 674 18163 800 18316
rect 866 18163 992 18316
rect 1058 18163 1184 18316
rect 1250 18163 1376 18316
rect 1828 18163 1860 18316
rect 1926 18163 2052 18316
rect 2118 18163 2244 18316
rect 2310 18163 2436 18316
rect 2502 18163 2628 18316
rect 2694 18163 2820 18316
rect 2886 18163 3012 18316
rect 3078 18163 3204 18316
rect 3656 18163 3688 18316
rect 3754 18163 3880 18316
rect 3946 18163 4072 18316
rect 4138 18163 4264 18316
rect 4330 18163 4456 18316
rect 4522 18163 4648 18316
rect 4714 18163 4840 18316
rect 4906 18163 5032 18316
rect 5484 18163 5516 18316
rect 5582 18163 5708 18316
rect 5774 18163 5900 18316
rect 5966 18163 6092 18316
rect 6158 18163 6284 18316
rect 6350 18163 6476 18316
rect 6542 18163 6668 18316
rect 6734 18163 6860 18316
rect 7312 18163 7344 18316
rect 7410 18163 7536 18316
rect 7602 18163 7728 18316
rect 7794 18163 7920 18316
rect 7986 18163 8112 18316
rect 8178 18163 8304 18316
rect 8370 18163 8496 18316
rect 8562 18163 8688 18316
rect 9140 18163 9172 18316
rect 9238 18163 9364 18316
rect 9430 18163 9556 18316
rect 9622 18163 9748 18316
rect 9814 18163 9940 18316
rect 10006 18163 10132 18316
rect 10198 18163 10324 18316
rect 10390 18163 10516 18316
rect 10968 18163 11000 18316
rect 11066 18163 11192 18316
rect 11258 18163 11384 18316
rect 11450 18163 11576 18316
rect 11642 18163 11768 18316
rect 11834 18163 11960 18316
rect 12026 18163 12152 18316
rect 12218 18163 12344 18316
rect 12796 18163 12828 18316
rect 12894 18163 13020 18316
rect 13086 18163 13212 18316
rect 13278 18163 13404 18316
rect 13470 18163 13596 18316
rect 13662 18163 13788 18316
rect 13854 18163 13980 18316
rect 14046 18163 14172 18316
rect 14624 18163 14656 18316
rect 14722 18163 14848 18316
rect 14914 18163 15040 18316
rect 15106 18163 15232 18316
rect 15298 18163 15424 18316
rect 15490 18163 15616 18316
rect 15682 18163 15808 18316
rect 15874 18163 16000 18316
rect 16452 18163 16484 18316
rect 16550 18163 16676 18316
rect 16742 18163 16868 18316
rect 16934 18163 17060 18316
rect 17126 18163 17252 18316
rect 17318 18163 17444 18316
rect 17510 18163 17636 18316
rect 17702 18163 17828 18316
rect 18280 18163 18312 18316
rect 18378 18163 18504 18316
rect 18570 18163 18696 18316
rect 18762 18163 18888 18316
rect 18954 18163 19080 18316
rect 19146 18163 19272 18316
rect 19338 18163 19464 18316
rect 19530 18163 19656 18316
rect 20108 18163 20140 18316
rect 20206 18163 20332 18316
rect 20398 18163 20524 18316
rect 20590 18163 20716 18316
rect 20782 18163 20908 18316
rect 20974 18163 21100 18316
rect 21166 18163 21292 18316
rect 21358 18163 21484 18316
rect 32 18153 98 18163
rect 224 18153 290 18163
rect 416 18153 482 18163
rect 608 18153 674 18163
rect 800 18153 866 18163
rect 992 18153 1058 18163
rect 1184 18153 1250 18163
rect 1376 18153 1442 18163
rect 1860 18153 1926 18163
rect 2052 18153 2118 18163
rect 2244 18153 2310 18163
rect 2436 18153 2502 18163
rect 2628 18153 2694 18163
rect 2820 18153 2886 18163
rect 3012 18153 3078 18163
rect 3204 18153 3270 18163
rect 3688 18153 3754 18163
rect 3880 18153 3946 18163
rect 4072 18153 4138 18163
rect 4264 18153 4330 18163
rect 4456 18153 4522 18163
rect 4648 18153 4714 18163
rect 4840 18153 4906 18163
rect 5032 18153 5098 18163
rect 5516 18153 5582 18163
rect 5708 18153 5774 18163
rect 5900 18153 5966 18163
rect 6092 18153 6158 18163
rect 6284 18153 6350 18163
rect 6476 18153 6542 18163
rect 6668 18153 6734 18163
rect 6860 18153 6926 18163
rect 7344 18153 7410 18163
rect 7536 18153 7602 18163
rect 7728 18153 7794 18163
rect 7920 18153 7986 18163
rect 8112 18153 8178 18163
rect 8304 18153 8370 18163
rect 8496 18153 8562 18163
rect 8688 18153 8754 18163
rect 9172 18153 9238 18163
rect 9364 18153 9430 18163
rect 9556 18153 9622 18163
rect 9748 18153 9814 18163
rect 9940 18153 10006 18163
rect 10132 18153 10198 18163
rect 10324 18153 10390 18163
rect 10516 18153 10582 18163
rect 11000 18153 11066 18163
rect 11192 18153 11258 18163
rect 11384 18153 11450 18163
rect 11576 18153 11642 18163
rect 11768 18153 11834 18163
rect 11960 18153 12026 18163
rect 12152 18153 12218 18163
rect 12344 18153 12410 18163
rect 12828 18153 12894 18163
rect 13020 18153 13086 18163
rect 13212 18153 13278 18163
rect 13404 18153 13470 18163
rect 13596 18153 13662 18163
rect 13788 18153 13854 18163
rect 13980 18153 14046 18163
rect 14172 18153 14238 18163
rect 14656 18153 14722 18163
rect 14848 18153 14914 18163
rect 15040 18153 15106 18163
rect 15232 18153 15298 18163
rect 15424 18153 15490 18163
rect 15616 18153 15682 18163
rect 15808 18153 15874 18163
rect 16000 18153 16066 18163
rect 16484 18153 16550 18163
rect 16676 18153 16742 18163
rect 16868 18153 16934 18163
rect 17060 18153 17126 18163
rect 17252 18153 17318 18163
rect 17444 18153 17510 18163
rect 17636 18153 17702 18163
rect 17828 18153 17894 18163
rect 18312 18153 18378 18163
rect 18504 18153 18570 18163
rect 18696 18153 18762 18163
rect 18888 18153 18954 18163
rect 19080 18153 19146 18163
rect 19272 18153 19338 18163
rect 19464 18153 19530 18163
rect 19656 18153 19722 18163
rect 20140 18153 20206 18163
rect 20332 18153 20398 18163
rect 20524 18153 20590 18163
rect 20716 18153 20782 18163
rect 20908 18153 20974 18163
rect 21100 18153 21166 18163
rect 21292 18153 21358 18163
rect 21484 18153 21550 18163
rect 128 18103 194 18113
rect 320 18103 386 18113
rect 512 18103 578 18113
rect 704 18103 770 18113
rect 896 18103 962 18113
rect 1088 18103 1154 18113
rect 1280 18103 1346 18113
rect 1472 18103 1528 18113
rect 1956 18103 2022 18113
rect 2148 18103 2214 18113
rect 2340 18103 2406 18113
rect 2532 18103 2598 18113
rect 2724 18103 2790 18113
rect 2916 18103 2982 18113
rect 3108 18103 3174 18113
rect 3300 18103 3356 18113
rect 3784 18103 3850 18113
rect 3976 18103 4042 18113
rect 4168 18103 4234 18113
rect 4360 18103 4426 18113
rect 4552 18103 4618 18113
rect 4744 18103 4810 18113
rect 4936 18103 5002 18113
rect 5128 18103 5184 18113
rect 5612 18103 5678 18113
rect 5804 18103 5870 18113
rect 5996 18103 6062 18113
rect 6188 18103 6254 18113
rect 6380 18103 6446 18113
rect 6572 18103 6638 18113
rect 6764 18103 6830 18113
rect 6956 18103 7012 18113
rect 7440 18103 7506 18113
rect 7632 18103 7698 18113
rect 7824 18103 7890 18113
rect 8016 18103 8082 18113
rect 8208 18103 8274 18113
rect 8400 18103 8466 18113
rect 8592 18103 8658 18113
rect 8784 18103 8840 18113
rect 9268 18103 9334 18113
rect 9460 18103 9526 18113
rect 9652 18103 9718 18113
rect 9844 18103 9910 18113
rect 10036 18103 10102 18113
rect 10228 18103 10294 18113
rect 10420 18103 10486 18113
rect 10612 18103 10668 18113
rect 11096 18103 11162 18113
rect 11288 18103 11354 18113
rect 11480 18103 11546 18113
rect 11672 18103 11738 18113
rect 11864 18103 11930 18113
rect 12056 18103 12122 18113
rect 12248 18103 12314 18113
rect 12440 18103 12496 18113
rect 12924 18103 12990 18113
rect 13116 18103 13182 18113
rect 13308 18103 13374 18113
rect 13500 18103 13566 18113
rect 13692 18103 13758 18113
rect 13884 18103 13950 18113
rect 14076 18103 14142 18113
rect 14268 18103 14324 18113
rect 14752 18103 14818 18113
rect 14944 18103 15010 18113
rect 15136 18103 15202 18113
rect 15328 18103 15394 18113
rect 15520 18103 15586 18113
rect 15712 18103 15778 18113
rect 15904 18103 15970 18113
rect 16096 18103 16152 18113
rect 16580 18103 16646 18113
rect 16772 18103 16838 18113
rect 16964 18103 17030 18113
rect 17156 18103 17222 18113
rect 17348 18103 17414 18113
rect 17540 18103 17606 18113
rect 17732 18103 17798 18113
rect 17924 18103 17980 18113
rect 18408 18103 18474 18113
rect 18600 18103 18666 18113
rect 18792 18103 18858 18113
rect 18984 18103 19050 18113
rect 19176 18103 19242 18113
rect 19368 18103 19434 18113
rect 19560 18103 19626 18113
rect 19752 18103 19808 18113
rect 20236 18103 20302 18113
rect 20428 18103 20494 18113
rect 20620 18103 20686 18113
rect 20812 18103 20878 18113
rect 21004 18103 21070 18113
rect 21196 18103 21262 18113
rect 21388 18103 21454 18113
rect 21580 18103 21636 18113
rect 0 17950 128 18103
rect 194 17950 320 18103
rect 386 17950 512 18103
rect 578 17950 704 18103
rect 770 17950 896 18103
rect 962 17950 1088 18103
rect 1154 17950 1280 18103
rect 1346 17950 1472 18103
rect 1528 17950 1708 18103
rect 1828 17950 1956 18103
rect 2022 17950 2148 18103
rect 2214 17950 2340 18103
rect 2406 17950 2532 18103
rect 2598 17950 2724 18103
rect 2790 17950 2916 18103
rect 2982 17950 3108 18103
rect 3174 17950 3300 18103
rect 3356 17950 3536 18103
rect 3656 17950 3784 18103
rect 3850 17950 3976 18103
rect 4042 17950 4168 18103
rect 4234 17950 4360 18103
rect 4426 17950 4552 18103
rect 4618 17950 4744 18103
rect 4810 17950 4936 18103
rect 5002 17950 5128 18103
rect 5184 17950 5364 18103
rect 5484 17950 5612 18103
rect 5678 17950 5804 18103
rect 5870 17950 5996 18103
rect 6062 17950 6188 18103
rect 6254 17950 6380 18103
rect 6446 17950 6572 18103
rect 6638 17950 6764 18103
rect 6830 17950 6956 18103
rect 7012 17950 7192 18103
rect 7312 17950 7440 18103
rect 7506 17950 7632 18103
rect 7698 17950 7824 18103
rect 7890 17950 8016 18103
rect 8082 17950 8208 18103
rect 8274 17950 8400 18103
rect 8466 17950 8592 18103
rect 8658 17950 8784 18103
rect 8840 17950 9020 18103
rect 9140 17950 9268 18103
rect 9334 17950 9460 18103
rect 9526 17950 9652 18103
rect 9718 17950 9844 18103
rect 9910 17950 10036 18103
rect 10102 17950 10228 18103
rect 10294 17950 10420 18103
rect 10486 17950 10612 18103
rect 10668 17950 10848 18103
rect 10968 17950 11096 18103
rect 11162 17950 11288 18103
rect 11354 17950 11480 18103
rect 11546 17950 11672 18103
rect 11738 17950 11864 18103
rect 11930 17950 12056 18103
rect 12122 17950 12248 18103
rect 12314 17950 12440 18103
rect 12496 17950 12676 18103
rect 12796 17950 12924 18103
rect 12990 17950 13116 18103
rect 13182 17950 13308 18103
rect 13374 17950 13500 18103
rect 13566 17950 13692 18103
rect 13758 17950 13884 18103
rect 13950 17950 14076 18103
rect 14142 17950 14268 18103
rect 14324 17950 14504 18103
rect 14624 17950 14752 18103
rect 14818 17950 14944 18103
rect 15010 17950 15136 18103
rect 15202 17950 15328 18103
rect 15394 17950 15520 18103
rect 15586 17950 15712 18103
rect 15778 17950 15904 18103
rect 15970 17950 16096 18103
rect 16152 17950 16332 18103
rect 16452 17950 16580 18103
rect 16646 17950 16772 18103
rect 16838 17950 16964 18103
rect 17030 17950 17156 18103
rect 17222 17950 17348 18103
rect 17414 17950 17540 18103
rect 17606 17950 17732 18103
rect 17798 17950 17924 18103
rect 17980 17950 18160 18103
rect 18280 17950 18408 18103
rect 18474 17950 18600 18103
rect 18666 17950 18792 18103
rect 18858 17950 18984 18103
rect 19050 17950 19176 18103
rect 19242 17950 19368 18103
rect 19434 17950 19560 18103
rect 19626 17950 19752 18103
rect 19808 17950 19988 18103
rect 20108 17950 20236 18103
rect 20302 17950 20428 18103
rect 20494 17950 20620 18103
rect 20686 17950 20812 18103
rect 20878 17950 21004 18103
rect 21070 17950 21196 18103
rect 21262 17950 21388 18103
rect 21454 17950 21580 18103
rect 21636 17950 21816 18103
rect 128 17940 194 17950
rect 320 17940 386 17950
rect 512 17940 578 17950
rect 704 17940 770 17950
rect 896 17940 962 17950
rect 1088 17940 1154 17950
rect 1280 17940 1346 17950
rect 1472 17940 1528 17950
rect 1956 17940 2022 17950
rect 2148 17940 2214 17950
rect 2340 17940 2406 17950
rect 2532 17940 2598 17950
rect 2724 17940 2790 17950
rect 2916 17940 2982 17950
rect 3108 17940 3174 17950
rect 3300 17940 3356 17950
rect 3784 17940 3850 17950
rect 3976 17940 4042 17950
rect 4168 17940 4234 17950
rect 4360 17940 4426 17950
rect 4552 17940 4618 17950
rect 4744 17940 4810 17950
rect 4936 17940 5002 17950
rect 5128 17940 5184 17950
rect 5612 17940 5678 17950
rect 5804 17940 5870 17950
rect 5996 17940 6062 17950
rect 6188 17940 6254 17950
rect 6380 17940 6446 17950
rect 6572 17940 6638 17950
rect 6764 17940 6830 17950
rect 6956 17940 7012 17950
rect 7440 17940 7506 17950
rect 7632 17940 7698 17950
rect 7824 17940 7890 17950
rect 8016 17940 8082 17950
rect 8208 17940 8274 17950
rect 8400 17940 8466 17950
rect 8592 17940 8658 17950
rect 8784 17940 8840 17950
rect 9268 17940 9334 17950
rect 9460 17940 9526 17950
rect 9652 17940 9718 17950
rect 9844 17940 9910 17950
rect 10036 17940 10102 17950
rect 10228 17940 10294 17950
rect 10420 17940 10486 17950
rect 10612 17940 10668 17950
rect 11096 17940 11162 17950
rect 11288 17940 11354 17950
rect 11480 17940 11546 17950
rect 11672 17940 11738 17950
rect 11864 17940 11930 17950
rect 12056 17940 12122 17950
rect 12248 17940 12314 17950
rect 12440 17940 12496 17950
rect 12924 17940 12990 17950
rect 13116 17940 13182 17950
rect 13308 17940 13374 17950
rect 13500 17940 13566 17950
rect 13692 17940 13758 17950
rect 13884 17940 13950 17950
rect 14076 17940 14142 17950
rect 14268 17940 14324 17950
rect 14752 17940 14818 17950
rect 14944 17940 15010 17950
rect 15136 17940 15202 17950
rect 15328 17940 15394 17950
rect 15520 17940 15586 17950
rect 15712 17940 15778 17950
rect 15904 17940 15970 17950
rect 16096 17940 16152 17950
rect 16580 17940 16646 17950
rect 16772 17940 16838 17950
rect 16964 17940 17030 17950
rect 17156 17940 17222 17950
rect 17348 17940 17414 17950
rect 17540 17940 17606 17950
rect 17732 17940 17798 17950
rect 17924 17940 17980 17950
rect 18408 17940 18474 17950
rect 18600 17940 18666 17950
rect 18792 17940 18858 17950
rect 18984 17940 19050 17950
rect 19176 17940 19242 17950
rect 19368 17940 19434 17950
rect 19560 17940 19626 17950
rect 19752 17940 19808 17950
rect 20236 17940 20302 17950
rect 20428 17940 20494 17950
rect 20620 17940 20686 17950
rect 20812 17940 20878 17950
rect 21004 17940 21070 17950
rect 21196 17940 21262 17950
rect 21388 17940 21454 17950
rect 21580 17940 21636 17950
rect 32 17602 98 17612
rect 224 17602 290 17612
rect 416 17602 482 17612
rect 608 17602 674 17612
rect 800 17602 866 17612
rect 992 17602 1058 17612
rect 1184 17602 1250 17612
rect 1376 17602 1442 17612
rect 1860 17602 1926 17612
rect 2052 17602 2118 17612
rect 2244 17602 2310 17612
rect 2436 17602 2502 17612
rect 2628 17602 2694 17612
rect 2820 17602 2886 17612
rect 3012 17602 3078 17612
rect 3204 17602 3270 17612
rect 3688 17602 3754 17612
rect 3880 17602 3946 17612
rect 4072 17602 4138 17612
rect 4264 17602 4330 17612
rect 4456 17602 4522 17612
rect 4648 17602 4714 17612
rect 4840 17602 4906 17612
rect 5032 17602 5098 17612
rect 5516 17602 5582 17612
rect 5708 17602 5774 17612
rect 5900 17602 5966 17612
rect 6092 17602 6158 17612
rect 6284 17602 6350 17612
rect 6476 17602 6542 17612
rect 6668 17602 6734 17612
rect 6860 17602 6926 17612
rect 7344 17602 7410 17612
rect 7536 17602 7602 17612
rect 7728 17602 7794 17612
rect 7920 17602 7986 17612
rect 8112 17602 8178 17612
rect 8304 17602 8370 17612
rect 8496 17602 8562 17612
rect 8688 17602 8754 17612
rect 9172 17602 9238 17612
rect 9364 17602 9430 17612
rect 9556 17602 9622 17612
rect 9748 17602 9814 17612
rect 9940 17602 10006 17612
rect 10132 17602 10198 17612
rect 10324 17602 10390 17612
rect 10516 17602 10582 17612
rect 11000 17602 11066 17612
rect 11192 17602 11258 17612
rect 11384 17602 11450 17612
rect 11576 17602 11642 17612
rect 11768 17602 11834 17612
rect 11960 17602 12026 17612
rect 12152 17602 12218 17612
rect 12344 17602 12410 17612
rect 12828 17602 12894 17612
rect 13020 17602 13086 17612
rect 13212 17602 13278 17612
rect 13404 17602 13470 17612
rect 13596 17602 13662 17612
rect 13788 17602 13854 17612
rect 13980 17602 14046 17612
rect 14172 17602 14238 17612
rect 14656 17602 14722 17612
rect 14848 17602 14914 17612
rect 15040 17602 15106 17612
rect 15232 17602 15298 17612
rect 15424 17602 15490 17612
rect 15616 17602 15682 17612
rect 15808 17602 15874 17612
rect 16000 17602 16066 17612
rect 16484 17602 16550 17612
rect 16676 17602 16742 17612
rect 16868 17602 16934 17612
rect 17060 17602 17126 17612
rect 17252 17602 17318 17612
rect 17444 17602 17510 17612
rect 17636 17602 17702 17612
rect 17828 17602 17894 17612
rect 18312 17602 18378 17612
rect 18504 17602 18570 17612
rect 18696 17602 18762 17612
rect 18888 17602 18954 17612
rect 19080 17602 19146 17612
rect 19272 17602 19338 17612
rect 19464 17602 19530 17612
rect 19656 17602 19722 17612
rect 20140 17602 20206 17612
rect 20332 17602 20398 17612
rect 20524 17602 20590 17612
rect 20716 17602 20782 17612
rect 20908 17602 20974 17612
rect 21100 17602 21166 17612
rect 21292 17602 21358 17612
rect 21484 17602 21550 17612
rect 0 17449 32 17602
rect 98 17449 224 17602
rect 290 17449 416 17602
rect 482 17449 608 17602
rect 674 17449 800 17602
rect 866 17449 992 17602
rect 1058 17449 1184 17602
rect 1250 17449 1376 17602
rect 1828 17449 1860 17602
rect 1926 17449 2052 17602
rect 2118 17449 2244 17602
rect 2310 17449 2436 17602
rect 2502 17449 2628 17602
rect 2694 17449 2820 17602
rect 2886 17449 3012 17602
rect 3078 17449 3204 17602
rect 3656 17449 3688 17602
rect 3754 17449 3880 17602
rect 3946 17449 4072 17602
rect 4138 17449 4264 17602
rect 4330 17449 4456 17602
rect 4522 17449 4648 17602
rect 4714 17449 4840 17602
rect 4906 17449 5032 17602
rect 5484 17449 5516 17602
rect 5582 17449 5708 17602
rect 5774 17449 5900 17602
rect 5966 17449 6092 17602
rect 6158 17449 6284 17602
rect 6350 17449 6476 17602
rect 6542 17449 6668 17602
rect 6734 17449 6860 17602
rect 7312 17449 7344 17602
rect 7410 17449 7536 17602
rect 7602 17449 7728 17602
rect 7794 17449 7920 17602
rect 7986 17449 8112 17602
rect 8178 17449 8304 17602
rect 8370 17449 8496 17602
rect 8562 17449 8688 17602
rect 9140 17449 9172 17602
rect 9238 17449 9364 17602
rect 9430 17449 9556 17602
rect 9622 17449 9748 17602
rect 9814 17449 9940 17602
rect 10006 17449 10132 17602
rect 10198 17449 10324 17602
rect 10390 17449 10516 17602
rect 10968 17449 11000 17602
rect 11066 17449 11192 17602
rect 11258 17449 11384 17602
rect 11450 17449 11576 17602
rect 11642 17449 11768 17602
rect 11834 17449 11960 17602
rect 12026 17449 12152 17602
rect 12218 17449 12344 17602
rect 12796 17449 12828 17602
rect 12894 17449 13020 17602
rect 13086 17449 13212 17602
rect 13278 17449 13404 17602
rect 13470 17449 13596 17602
rect 13662 17449 13788 17602
rect 13854 17449 13980 17602
rect 14046 17449 14172 17602
rect 14624 17449 14656 17602
rect 14722 17449 14848 17602
rect 14914 17449 15040 17602
rect 15106 17449 15232 17602
rect 15298 17449 15424 17602
rect 15490 17449 15616 17602
rect 15682 17449 15808 17602
rect 15874 17449 16000 17602
rect 16452 17449 16484 17602
rect 16550 17449 16676 17602
rect 16742 17449 16868 17602
rect 16934 17449 17060 17602
rect 17126 17449 17252 17602
rect 17318 17449 17444 17602
rect 17510 17449 17636 17602
rect 17702 17449 17828 17602
rect 18280 17449 18312 17602
rect 18378 17449 18504 17602
rect 18570 17449 18696 17602
rect 18762 17449 18888 17602
rect 18954 17449 19080 17602
rect 19146 17449 19272 17602
rect 19338 17449 19464 17602
rect 19530 17449 19656 17602
rect 20108 17449 20140 17602
rect 20206 17449 20332 17602
rect 20398 17449 20524 17602
rect 20590 17449 20716 17602
rect 20782 17449 20908 17602
rect 20974 17449 21100 17602
rect 21166 17449 21292 17602
rect 21358 17449 21484 17602
rect 32 17439 98 17449
rect 224 17439 290 17449
rect 416 17439 482 17449
rect 608 17439 674 17449
rect 800 17439 866 17449
rect 992 17439 1058 17449
rect 1184 17439 1250 17449
rect 1376 17439 1442 17449
rect 1860 17439 1926 17449
rect 2052 17439 2118 17449
rect 2244 17439 2310 17449
rect 2436 17439 2502 17449
rect 2628 17439 2694 17449
rect 2820 17439 2886 17449
rect 3012 17439 3078 17449
rect 3204 17439 3270 17449
rect 3688 17439 3754 17449
rect 3880 17439 3946 17449
rect 4072 17439 4138 17449
rect 4264 17439 4330 17449
rect 4456 17439 4522 17449
rect 4648 17439 4714 17449
rect 4840 17439 4906 17449
rect 5032 17439 5098 17449
rect 5516 17439 5582 17449
rect 5708 17439 5774 17449
rect 5900 17439 5966 17449
rect 6092 17439 6158 17449
rect 6284 17439 6350 17449
rect 6476 17439 6542 17449
rect 6668 17439 6734 17449
rect 6860 17439 6926 17449
rect 7344 17439 7410 17449
rect 7536 17439 7602 17449
rect 7728 17439 7794 17449
rect 7920 17439 7986 17449
rect 8112 17439 8178 17449
rect 8304 17439 8370 17449
rect 8496 17439 8562 17449
rect 8688 17439 8754 17449
rect 9172 17439 9238 17449
rect 9364 17439 9430 17449
rect 9556 17439 9622 17449
rect 9748 17439 9814 17449
rect 9940 17439 10006 17449
rect 10132 17439 10198 17449
rect 10324 17439 10390 17449
rect 10516 17439 10582 17449
rect 11000 17439 11066 17449
rect 11192 17439 11258 17449
rect 11384 17439 11450 17449
rect 11576 17439 11642 17449
rect 11768 17439 11834 17449
rect 11960 17439 12026 17449
rect 12152 17439 12218 17449
rect 12344 17439 12410 17449
rect 12828 17439 12894 17449
rect 13020 17439 13086 17449
rect 13212 17439 13278 17449
rect 13404 17439 13470 17449
rect 13596 17439 13662 17449
rect 13788 17439 13854 17449
rect 13980 17439 14046 17449
rect 14172 17439 14238 17449
rect 14656 17439 14722 17449
rect 14848 17439 14914 17449
rect 15040 17439 15106 17449
rect 15232 17439 15298 17449
rect 15424 17439 15490 17449
rect 15616 17439 15682 17449
rect 15808 17439 15874 17449
rect 16000 17439 16066 17449
rect 16484 17439 16550 17449
rect 16676 17439 16742 17449
rect 16868 17439 16934 17449
rect 17060 17439 17126 17449
rect 17252 17439 17318 17449
rect 17444 17439 17510 17449
rect 17636 17439 17702 17449
rect 17828 17439 17894 17449
rect 18312 17439 18378 17449
rect 18504 17439 18570 17449
rect 18696 17439 18762 17449
rect 18888 17439 18954 17449
rect 19080 17439 19146 17449
rect 19272 17439 19338 17449
rect 19464 17439 19530 17449
rect 19656 17439 19722 17449
rect 20140 17439 20206 17449
rect 20332 17439 20398 17449
rect 20524 17439 20590 17449
rect 20716 17439 20782 17449
rect 20908 17439 20974 17449
rect 21100 17439 21166 17449
rect 21292 17439 21358 17449
rect 21484 17439 21550 17449
rect 128 17389 194 17399
rect 320 17389 386 17399
rect 512 17389 578 17399
rect 704 17389 770 17399
rect 896 17389 962 17399
rect 1088 17389 1154 17399
rect 1280 17389 1346 17399
rect 1472 17389 1528 17399
rect 1956 17389 2022 17399
rect 2148 17389 2214 17399
rect 2340 17389 2406 17399
rect 2532 17389 2598 17399
rect 2724 17389 2790 17399
rect 2916 17389 2982 17399
rect 3108 17389 3174 17399
rect 3300 17389 3356 17399
rect 3784 17389 3850 17399
rect 3976 17389 4042 17399
rect 4168 17389 4234 17399
rect 4360 17389 4426 17399
rect 4552 17389 4618 17399
rect 4744 17389 4810 17399
rect 4936 17389 5002 17399
rect 5128 17389 5184 17399
rect 5612 17389 5678 17399
rect 5804 17389 5870 17399
rect 5996 17389 6062 17399
rect 6188 17389 6254 17399
rect 6380 17389 6446 17399
rect 6572 17389 6638 17399
rect 6764 17389 6830 17399
rect 6956 17389 7012 17399
rect 7440 17389 7506 17399
rect 7632 17389 7698 17399
rect 7824 17389 7890 17399
rect 8016 17389 8082 17399
rect 8208 17389 8274 17399
rect 8400 17389 8466 17399
rect 8592 17389 8658 17399
rect 8784 17389 8840 17399
rect 9268 17389 9334 17399
rect 9460 17389 9526 17399
rect 9652 17389 9718 17399
rect 9844 17389 9910 17399
rect 10036 17389 10102 17399
rect 10228 17389 10294 17399
rect 10420 17389 10486 17399
rect 10612 17389 10668 17399
rect 11096 17389 11162 17399
rect 11288 17389 11354 17399
rect 11480 17389 11546 17399
rect 11672 17389 11738 17399
rect 11864 17389 11930 17399
rect 12056 17389 12122 17399
rect 12248 17389 12314 17399
rect 12440 17389 12496 17399
rect 12924 17389 12990 17399
rect 13116 17389 13182 17399
rect 13308 17389 13374 17399
rect 13500 17389 13566 17399
rect 13692 17389 13758 17399
rect 13884 17389 13950 17399
rect 14076 17389 14142 17399
rect 14268 17389 14324 17399
rect 14752 17389 14818 17399
rect 14944 17389 15010 17399
rect 15136 17389 15202 17399
rect 15328 17389 15394 17399
rect 15520 17389 15586 17399
rect 15712 17389 15778 17399
rect 15904 17389 15970 17399
rect 16096 17389 16152 17399
rect 16580 17389 16646 17399
rect 16772 17389 16838 17399
rect 16964 17389 17030 17399
rect 17156 17389 17222 17399
rect 17348 17389 17414 17399
rect 17540 17389 17606 17399
rect 17732 17389 17798 17399
rect 17924 17389 17980 17399
rect 18408 17389 18474 17399
rect 18600 17389 18666 17399
rect 18792 17389 18858 17399
rect 18984 17389 19050 17399
rect 19176 17389 19242 17399
rect 19368 17389 19434 17399
rect 19560 17389 19626 17399
rect 19752 17389 19808 17399
rect 20236 17389 20302 17399
rect 20428 17389 20494 17399
rect 20620 17389 20686 17399
rect 20812 17389 20878 17399
rect 21004 17389 21070 17399
rect 21196 17389 21262 17399
rect 21388 17389 21454 17399
rect 21580 17389 21636 17399
rect 0 17236 128 17389
rect 194 17236 320 17389
rect 386 17236 512 17389
rect 578 17236 704 17389
rect 770 17236 896 17389
rect 962 17236 1088 17389
rect 1154 17236 1280 17389
rect 1346 17236 1472 17389
rect 1528 17236 1708 17389
rect 1828 17236 1956 17389
rect 2022 17236 2148 17389
rect 2214 17236 2340 17389
rect 2406 17236 2532 17389
rect 2598 17236 2724 17389
rect 2790 17236 2916 17389
rect 2982 17236 3108 17389
rect 3174 17236 3300 17389
rect 3356 17236 3536 17389
rect 3656 17236 3784 17389
rect 3850 17236 3976 17389
rect 4042 17236 4168 17389
rect 4234 17236 4360 17389
rect 4426 17236 4552 17389
rect 4618 17236 4744 17389
rect 4810 17236 4936 17389
rect 5002 17236 5128 17389
rect 5184 17236 5364 17389
rect 5484 17236 5612 17389
rect 5678 17236 5804 17389
rect 5870 17236 5996 17389
rect 6062 17236 6188 17389
rect 6254 17236 6380 17389
rect 6446 17236 6572 17389
rect 6638 17236 6764 17389
rect 6830 17236 6956 17389
rect 7012 17236 7192 17389
rect 7312 17236 7440 17389
rect 7506 17236 7632 17389
rect 7698 17236 7824 17389
rect 7890 17236 8016 17389
rect 8082 17236 8208 17389
rect 8274 17236 8400 17389
rect 8466 17236 8592 17389
rect 8658 17236 8784 17389
rect 8840 17236 9020 17389
rect 9140 17236 9268 17389
rect 9334 17236 9460 17389
rect 9526 17236 9652 17389
rect 9718 17236 9844 17389
rect 9910 17236 10036 17389
rect 10102 17236 10228 17389
rect 10294 17236 10420 17389
rect 10486 17236 10612 17389
rect 10668 17236 10848 17389
rect 10968 17236 11096 17389
rect 11162 17236 11288 17389
rect 11354 17236 11480 17389
rect 11546 17236 11672 17389
rect 11738 17236 11864 17389
rect 11930 17236 12056 17389
rect 12122 17236 12248 17389
rect 12314 17236 12440 17389
rect 12496 17236 12676 17389
rect 12796 17236 12924 17389
rect 12990 17236 13116 17389
rect 13182 17236 13308 17389
rect 13374 17236 13500 17389
rect 13566 17236 13692 17389
rect 13758 17236 13884 17389
rect 13950 17236 14076 17389
rect 14142 17236 14268 17389
rect 14324 17236 14504 17389
rect 14624 17236 14752 17389
rect 14818 17236 14944 17389
rect 15010 17236 15136 17389
rect 15202 17236 15328 17389
rect 15394 17236 15520 17389
rect 15586 17236 15712 17389
rect 15778 17236 15904 17389
rect 15970 17236 16096 17389
rect 16152 17236 16332 17389
rect 16452 17236 16580 17389
rect 16646 17236 16772 17389
rect 16838 17236 16964 17389
rect 17030 17236 17156 17389
rect 17222 17236 17348 17389
rect 17414 17236 17540 17389
rect 17606 17236 17732 17389
rect 17798 17236 17924 17389
rect 17980 17236 18160 17389
rect 18280 17236 18408 17389
rect 18474 17236 18600 17389
rect 18666 17236 18792 17389
rect 18858 17236 18984 17389
rect 19050 17236 19176 17389
rect 19242 17236 19368 17389
rect 19434 17236 19560 17389
rect 19626 17236 19752 17389
rect 19808 17236 19988 17389
rect 20108 17236 20236 17389
rect 20302 17236 20428 17389
rect 20494 17236 20620 17389
rect 20686 17236 20812 17389
rect 20878 17236 21004 17389
rect 21070 17236 21196 17389
rect 21262 17236 21388 17389
rect 21454 17236 21580 17389
rect 21636 17236 21816 17389
rect 128 17226 194 17236
rect 320 17226 386 17236
rect 512 17226 578 17236
rect 704 17226 770 17236
rect 896 17226 962 17236
rect 1088 17226 1154 17236
rect 1280 17226 1346 17236
rect 1472 17226 1528 17236
rect 1956 17226 2022 17236
rect 2148 17226 2214 17236
rect 2340 17226 2406 17236
rect 2532 17226 2598 17236
rect 2724 17226 2790 17236
rect 2916 17226 2982 17236
rect 3108 17226 3174 17236
rect 3300 17226 3356 17236
rect 3784 17226 3850 17236
rect 3976 17226 4042 17236
rect 4168 17226 4234 17236
rect 4360 17226 4426 17236
rect 4552 17226 4618 17236
rect 4744 17226 4810 17236
rect 4936 17226 5002 17236
rect 5128 17226 5184 17236
rect 5612 17226 5678 17236
rect 5804 17226 5870 17236
rect 5996 17226 6062 17236
rect 6188 17226 6254 17236
rect 6380 17226 6446 17236
rect 6572 17226 6638 17236
rect 6764 17226 6830 17236
rect 6956 17226 7012 17236
rect 7440 17226 7506 17236
rect 7632 17226 7698 17236
rect 7824 17226 7890 17236
rect 8016 17226 8082 17236
rect 8208 17226 8274 17236
rect 8400 17226 8466 17236
rect 8592 17226 8658 17236
rect 8784 17226 8840 17236
rect 9268 17226 9334 17236
rect 9460 17226 9526 17236
rect 9652 17226 9718 17236
rect 9844 17226 9910 17236
rect 10036 17226 10102 17236
rect 10228 17226 10294 17236
rect 10420 17226 10486 17236
rect 10612 17226 10668 17236
rect 11096 17226 11162 17236
rect 11288 17226 11354 17236
rect 11480 17226 11546 17236
rect 11672 17226 11738 17236
rect 11864 17226 11930 17236
rect 12056 17226 12122 17236
rect 12248 17226 12314 17236
rect 12440 17226 12496 17236
rect 12924 17226 12990 17236
rect 13116 17226 13182 17236
rect 13308 17226 13374 17236
rect 13500 17226 13566 17236
rect 13692 17226 13758 17236
rect 13884 17226 13950 17236
rect 14076 17226 14142 17236
rect 14268 17226 14324 17236
rect 14752 17226 14818 17236
rect 14944 17226 15010 17236
rect 15136 17226 15202 17236
rect 15328 17226 15394 17236
rect 15520 17226 15586 17236
rect 15712 17226 15778 17236
rect 15904 17226 15970 17236
rect 16096 17226 16152 17236
rect 16580 17226 16646 17236
rect 16772 17226 16838 17236
rect 16964 17226 17030 17236
rect 17156 17226 17222 17236
rect 17348 17226 17414 17236
rect 17540 17226 17606 17236
rect 17732 17226 17798 17236
rect 17924 17226 17980 17236
rect 18408 17226 18474 17236
rect 18600 17226 18666 17236
rect 18792 17226 18858 17236
rect 18984 17226 19050 17236
rect 19176 17226 19242 17236
rect 19368 17226 19434 17236
rect 19560 17226 19626 17236
rect 19752 17226 19808 17236
rect 20236 17226 20302 17236
rect 20428 17226 20494 17236
rect 20620 17226 20686 17236
rect 20812 17226 20878 17236
rect 21004 17226 21070 17236
rect 21196 17226 21262 17236
rect 21388 17226 21454 17236
rect 21580 17226 21636 17236
rect 32 16888 98 16898
rect 224 16888 290 16898
rect 416 16888 482 16898
rect 608 16888 674 16898
rect 800 16888 866 16898
rect 992 16888 1058 16898
rect 1184 16888 1250 16898
rect 1376 16888 1442 16898
rect 1860 16888 1926 16898
rect 2052 16888 2118 16898
rect 2244 16888 2310 16898
rect 2436 16888 2502 16898
rect 2628 16888 2694 16898
rect 2820 16888 2886 16898
rect 3012 16888 3078 16898
rect 3204 16888 3270 16898
rect 3688 16888 3754 16898
rect 3880 16888 3946 16898
rect 4072 16888 4138 16898
rect 4264 16888 4330 16898
rect 4456 16888 4522 16898
rect 4648 16888 4714 16898
rect 4840 16888 4906 16898
rect 5032 16888 5098 16898
rect 5516 16888 5582 16898
rect 5708 16888 5774 16898
rect 5900 16888 5966 16898
rect 6092 16888 6158 16898
rect 6284 16888 6350 16898
rect 6476 16888 6542 16898
rect 6668 16888 6734 16898
rect 6860 16888 6926 16898
rect 7344 16888 7410 16898
rect 7536 16888 7602 16898
rect 7728 16888 7794 16898
rect 7920 16888 7986 16898
rect 8112 16888 8178 16898
rect 8304 16888 8370 16898
rect 8496 16888 8562 16898
rect 8688 16888 8754 16898
rect 9172 16888 9238 16898
rect 9364 16888 9430 16898
rect 9556 16888 9622 16898
rect 9748 16888 9814 16898
rect 9940 16888 10006 16898
rect 10132 16888 10198 16898
rect 10324 16888 10390 16898
rect 10516 16888 10582 16898
rect 11000 16888 11066 16898
rect 11192 16888 11258 16898
rect 11384 16888 11450 16898
rect 11576 16888 11642 16898
rect 11768 16888 11834 16898
rect 11960 16888 12026 16898
rect 12152 16888 12218 16898
rect 12344 16888 12410 16898
rect 12828 16888 12894 16898
rect 13020 16888 13086 16898
rect 13212 16888 13278 16898
rect 13404 16888 13470 16898
rect 13596 16888 13662 16898
rect 13788 16888 13854 16898
rect 13980 16888 14046 16898
rect 14172 16888 14238 16898
rect 14656 16888 14722 16898
rect 14848 16888 14914 16898
rect 15040 16888 15106 16898
rect 15232 16888 15298 16898
rect 15424 16888 15490 16898
rect 15616 16888 15682 16898
rect 15808 16888 15874 16898
rect 16000 16888 16066 16898
rect 16484 16888 16550 16898
rect 16676 16888 16742 16898
rect 16868 16888 16934 16898
rect 17060 16888 17126 16898
rect 17252 16888 17318 16898
rect 17444 16888 17510 16898
rect 17636 16888 17702 16898
rect 17828 16888 17894 16898
rect 18312 16888 18378 16898
rect 18504 16888 18570 16898
rect 18696 16888 18762 16898
rect 18888 16888 18954 16898
rect 19080 16888 19146 16898
rect 19272 16888 19338 16898
rect 19464 16888 19530 16898
rect 19656 16888 19722 16898
rect 20140 16888 20206 16898
rect 20332 16888 20398 16898
rect 20524 16888 20590 16898
rect 20716 16888 20782 16898
rect 20908 16888 20974 16898
rect 21100 16888 21166 16898
rect 21292 16888 21358 16898
rect 21484 16888 21550 16898
rect 0 16735 32 16888
rect 98 16735 224 16888
rect 290 16735 416 16888
rect 482 16735 608 16888
rect 674 16735 800 16888
rect 866 16735 992 16888
rect 1058 16735 1184 16888
rect 1250 16735 1376 16888
rect 1828 16735 1860 16888
rect 1926 16735 2052 16888
rect 2118 16735 2244 16888
rect 2310 16735 2436 16888
rect 2502 16735 2628 16888
rect 2694 16735 2820 16888
rect 2886 16735 3012 16888
rect 3078 16735 3204 16888
rect 3656 16735 3688 16888
rect 3754 16735 3880 16888
rect 3946 16735 4072 16888
rect 4138 16735 4264 16888
rect 4330 16735 4456 16888
rect 4522 16735 4648 16888
rect 4714 16735 4840 16888
rect 4906 16735 5032 16888
rect 5484 16735 5516 16888
rect 5582 16735 5708 16888
rect 5774 16735 5900 16888
rect 5966 16735 6092 16888
rect 6158 16735 6284 16888
rect 6350 16735 6476 16888
rect 6542 16735 6668 16888
rect 6734 16735 6860 16888
rect 7312 16735 7344 16888
rect 7410 16735 7536 16888
rect 7602 16735 7728 16888
rect 7794 16735 7920 16888
rect 7986 16735 8112 16888
rect 8178 16735 8304 16888
rect 8370 16735 8496 16888
rect 8562 16735 8688 16888
rect 9140 16735 9172 16888
rect 9238 16735 9364 16888
rect 9430 16735 9556 16888
rect 9622 16735 9748 16888
rect 9814 16735 9940 16888
rect 10006 16735 10132 16888
rect 10198 16735 10324 16888
rect 10390 16735 10516 16888
rect 10968 16735 11000 16888
rect 11066 16735 11192 16888
rect 11258 16735 11384 16888
rect 11450 16735 11576 16888
rect 11642 16735 11768 16888
rect 11834 16735 11960 16888
rect 12026 16735 12152 16888
rect 12218 16735 12344 16888
rect 12796 16735 12828 16888
rect 12894 16735 13020 16888
rect 13086 16735 13212 16888
rect 13278 16735 13404 16888
rect 13470 16735 13596 16888
rect 13662 16735 13788 16888
rect 13854 16735 13980 16888
rect 14046 16735 14172 16888
rect 14624 16735 14656 16888
rect 14722 16735 14848 16888
rect 14914 16735 15040 16888
rect 15106 16735 15232 16888
rect 15298 16735 15424 16888
rect 15490 16735 15616 16888
rect 15682 16735 15808 16888
rect 15874 16735 16000 16888
rect 16452 16735 16484 16888
rect 16550 16735 16676 16888
rect 16742 16735 16868 16888
rect 16934 16735 17060 16888
rect 17126 16735 17252 16888
rect 17318 16735 17444 16888
rect 17510 16735 17636 16888
rect 17702 16735 17828 16888
rect 18280 16735 18312 16888
rect 18378 16735 18504 16888
rect 18570 16735 18696 16888
rect 18762 16735 18888 16888
rect 18954 16735 19080 16888
rect 19146 16735 19272 16888
rect 19338 16735 19464 16888
rect 19530 16735 19656 16888
rect 20108 16735 20140 16888
rect 20206 16735 20332 16888
rect 20398 16735 20524 16888
rect 20590 16735 20716 16888
rect 20782 16735 20908 16888
rect 20974 16735 21100 16888
rect 21166 16735 21292 16888
rect 21358 16735 21484 16888
rect 32 16725 98 16735
rect 224 16725 290 16735
rect 416 16725 482 16735
rect 608 16725 674 16735
rect 800 16725 866 16735
rect 992 16725 1058 16735
rect 1184 16725 1250 16735
rect 1376 16725 1442 16735
rect 1860 16725 1926 16735
rect 2052 16725 2118 16735
rect 2244 16725 2310 16735
rect 2436 16725 2502 16735
rect 2628 16725 2694 16735
rect 2820 16725 2886 16735
rect 3012 16725 3078 16735
rect 3204 16725 3270 16735
rect 3688 16725 3754 16735
rect 3880 16725 3946 16735
rect 4072 16725 4138 16735
rect 4264 16725 4330 16735
rect 4456 16725 4522 16735
rect 4648 16725 4714 16735
rect 4840 16725 4906 16735
rect 5032 16725 5098 16735
rect 5516 16725 5582 16735
rect 5708 16725 5774 16735
rect 5900 16725 5966 16735
rect 6092 16725 6158 16735
rect 6284 16725 6350 16735
rect 6476 16725 6542 16735
rect 6668 16725 6734 16735
rect 6860 16725 6926 16735
rect 7344 16725 7410 16735
rect 7536 16725 7602 16735
rect 7728 16725 7794 16735
rect 7920 16725 7986 16735
rect 8112 16725 8178 16735
rect 8304 16725 8370 16735
rect 8496 16725 8562 16735
rect 8688 16725 8754 16735
rect 9172 16725 9238 16735
rect 9364 16725 9430 16735
rect 9556 16725 9622 16735
rect 9748 16725 9814 16735
rect 9940 16725 10006 16735
rect 10132 16725 10198 16735
rect 10324 16725 10390 16735
rect 10516 16725 10582 16735
rect 11000 16725 11066 16735
rect 11192 16725 11258 16735
rect 11384 16725 11450 16735
rect 11576 16725 11642 16735
rect 11768 16725 11834 16735
rect 11960 16725 12026 16735
rect 12152 16725 12218 16735
rect 12344 16725 12410 16735
rect 12828 16725 12894 16735
rect 13020 16725 13086 16735
rect 13212 16725 13278 16735
rect 13404 16725 13470 16735
rect 13596 16725 13662 16735
rect 13788 16725 13854 16735
rect 13980 16725 14046 16735
rect 14172 16725 14238 16735
rect 14656 16725 14722 16735
rect 14848 16725 14914 16735
rect 15040 16725 15106 16735
rect 15232 16725 15298 16735
rect 15424 16725 15490 16735
rect 15616 16725 15682 16735
rect 15808 16725 15874 16735
rect 16000 16725 16066 16735
rect 16484 16725 16550 16735
rect 16676 16725 16742 16735
rect 16868 16725 16934 16735
rect 17060 16725 17126 16735
rect 17252 16725 17318 16735
rect 17444 16725 17510 16735
rect 17636 16725 17702 16735
rect 17828 16725 17894 16735
rect 18312 16725 18378 16735
rect 18504 16725 18570 16735
rect 18696 16725 18762 16735
rect 18888 16725 18954 16735
rect 19080 16725 19146 16735
rect 19272 16725 19338 16735
rect 19464 16725 19530 16735
rect 19656 16725 19722 16735
rect 20140 16725 20206 16735
rect 20332 16725 20398 16735
rect 20524 16725 20590 16735
rect 20716 16725 20782 16735
rect 20908 16725 20974 16735
rect 21100 16725 21166 16735
rect 21292 16725 21358 16735
rect 21484 16725 21550 16735
rect 128 16675 194 16685
rect 320 16675 386 16685
rect 512 16675 578 16685
rect 704 16675 770 16685
rect 896 16675 962 16685
rect 1088 16675 1154 16685
rect 1280 16675 1346 16685
rect 1472 16675 1528 16685
rect 1956 16675 2022 16685
rect 2148 16675 2214 16685
rect 2340 16675 2406 16685
rect 2532 16675 2598 16685
rect 2724 16675 2790 16685
rect 2916 16675 2982 16685
rect 3108 16675 3174 16685
rect 3300 16675 3356 16685
rect 3784 16675 3850 16685
rect 3976 16675 4042 16685
rect 4168 16675 4234 16685
rect 4360 16675 4426 16685
rect 4552 16675 4618 16685
rect 4744 16675 4810 16685
rect 4936 16675 5002 16685
rect 5128 16675 5184 16685
rect 5612 16675 5678 16685
rect 5804 16675 5870 16685
rect 5996 16675 6062 16685
rect 6188 16675 6254 16685
rect 6380 16675 6446 16685
rect 6572 16675 6638 16685
rect 6764 16675 6830 16685
rect 6956 16675 7012 16685
rect 7440 16675 7506 16685
rect 7632 16675 7698 16685
rect 7824 16675 7890 16685
rect 8016 16675 8082 16685
rect 8208 16675 8274 16685
rect 8400 16675 8466 16685
rect 8592 16675 8658 16685
rect 8784 16675 8840 16685
rect 9268 16675 9334 16685
rect 9460 16675 9526 16685
rect 9652 16675 9718 16685
rect 9844 16675 9910 16685
rect 10036 16675 10102 16685
rect 10228 16675 10294 16685
rect 10420 16675 10486 16685
rect 10612 16675 10668 16685
rect 11096 16675 11162 16685
rect 11288 16675 11354 16685
rect 11480 16675 11546 16685
rect 11672 16675 11738 16685
rect 11864 16675 11930 16685
rect 12056 16675 12122 16685
rect 12248 16675 12314 16685
rect 12440 16675 12496 16685
rect 12924 16675 12990 16685
rect 13116 16675 13182 16685
rect 13308 16675 13374 16685
rect 13500 16675 13566 16685
rect 13692 16675 13758 16685
rect 13884 16675 13950 16685
rect 14076 16675 14142 16685
rect 14268 16675 14324 16685
rect 14752 16675 14818 16685
rect 14944 16675 15010 16685
rect 15136 16675 15202 16685
rect 15328 16675 15394 16685
rect 15520 16675 15586 16685
rect 15712 16675 15778 16685
rect 15904 16675 15970 16685
rect 16096 16675 16152 16685
rect 16580 16675 16646 16685
rect 16772 16675 16838 16685
rect 16964 16675 17030 16685
rect 17156 16675 17222 16685
rect 17348 16675 17414 16685
rect 17540 16675 17606 16685
rect 17732 16675 17798 16685
rect 17924 16675 17980 16685
rect 18408 16675 18474 16685
rect 18600 16675 18666 16685
rect 18792 16675 18858 16685
rect 18984 16675 19050 16685
rect 19176 16675 19242 16685
rect 19368 16675 19434 16685
rect 19560 16675 19626 16685
rect 19752 16675 19808 16685
rect 20236 16675 20302 16685
rect 20428 16675 20494 16685
rect 20620 16675 20686 16685
rect 20812 16675 20878 16685
rect 21004 16675 21070 16685
rect 21196 16675 21262 16685
rect 21388 16675 21454 16685
rect 21580 16675 21636 16685
rect 0 16522 128 16675
rect 194 16522 320 16675
rect 386 16522 512 16675
rect 578 16522 704 16675
rect 770 16522 896 16675
rect 962 16522 1088 16675
rect 1154 16522 1280 16675
rect 1346 16522 1472 16675
rect 1528 16522 1708 16675
rect 1828 16522 1956 16675
rect 2022 16522 2148 16675
rect 2214 16522 2340 16675
rect 2406 16522 2532 16675
rect 2598 16522 2724 16675
rect 2790 16522 2916 16675
rect 2982 16522 3108 16675
rect 3174 16522 3300 16675
rect 3356 16522 3536 16675
rect 3656 16522 3784 16675
rect 3850 16522 3976 16675
rect 4042 16522 4168 16675
rect 4234 16522 4360 16675
rect 4426 16522 4552 16675
rect 4618 16522 4744 16675
rect 4810 16522 4936 16675
rect 5002 16522 5128 16675
rect 5184 16522 5364 16675
rect 5484 16522 5612 16675
rect 5678 16522 5804 16675
rect 5870 16522 5996 16675
rect 6062 16522 6188 16675
rect 6254 16522 6380 16675
rect 6446 16522 6572 16675
rect 6638 16522 6764 16675
rect 6830 16522 6956 16675
rect 7012 16522 7192 16675
rect 7312 16522 7440 16675
rect 7506 16522 7632 16675
rect 7698 16522 7824 16675
rect 7890 16522 8016 16675
rect 8082 16522 8208 16675
rect 8274 16522 8400 16675
rect 8466 16522 8592 16675
rect 8658 16522 8784 16675
rect 8840 16522 9020 16675
rect 9140 16522 9268 16675
rect 9334 16522 9460 16675
rect 9526 16522 9652 16675
rect 9718 16522 9844 16675
rect 9910 16522 10036 16675
rect 10102 16522 10228 16675
rect 10294 16522 10420 16675
rect 10486 16522 10612 16675
rect 10668 16522 10848 16675
rect 10968 16522 11096 16675
rect 11162 16522 11288 16675
rect 11354 16522 11480 16675
rect 11546 16522 11672 16675
rect 11738 16522 11864 16675
rect 11930 16522 12056 16675
rect 12122 16522 12248 16675
rect 12314 16522 12440 16675
rect 12496 16522 12676 16675
rect 12796 16522 12924 16675
rect 12990 16522 13116 16675
rect 13182 16522 13308 16675
rect 13374 16522 13500 16675
rect 13566 16522 13692 16675
rect 13758 16522 13884 16675
rect 13950 16522 14076 16675
rect 14142 16522 14268 16675
rect 14324 16522 14504 16675
rect 14624 16522 14752 16675
rect 14818 16522 14944 16675
rect 15010 16522 15136 16675
rect 15202 16522 15328 16675
rect 15394 16522 15520 16675
rect 15586 16522 15712 16675
rect 15778 16522 15904 16675
rect 15970 16522 16096 16675
rect 16152 16522 16332 16675
rect 16452 16522 16580 16675
rect 16646 16522 16772 16675
rect 16838 16522 16964 16675
rect 17030 16522 17156 16675
rect 17222 16522 17348 16675
rect 17414 16522 17540 16675
rect 17606 16522 17732 16675
rect 17798 16522 17924 16675
rect 17980 16522 18160 16675
rect 18280 16522 18408 16675
rect 18474 16522 18600 16675
rect 18666 16522 18792 16675
rect 18858 16522 18984 16675
rect 19050 16522 19176 16675
rect 19242 16522 19368 16675
rect 19434 16522 19560 16675
rect 19626 16522 19752 16675
rect 19808 16522 19988 16675
rect 20108 16522 20236 16675
rect 20302 16522 20428 16675
rect 20494 16522 20620 16675
rect 20686 16522 20812 16675
rect 20878 16522 21004 16675
rect 21070 16522 21196 16675
rect 21262 16522 21388 16675
rect 21454 16522 21580 16675
rect 21636 16522 21816 16675
rect 128 16512 194 16522
rect 320 16512 386 16522
rect 512 16512 578 16522
rect 704 16512 770 16522
rect 896 16512 962 16522
rect 1088 16512 1154 16522
rect 1280 16512 1346 16522
rect 1472 16512 1528 16522
rect 1956 16512 2022 16522
rect 2148 16512 2214 16522
rect 2340 16512 2406 16522
rect 2532 16512 2598 16522
rect 2724 16512 2790 16522
rect 2916 16512 2982 16522
rect 3108 16512 3174 16522
rect 3300 16512 3356 16522
rect 3784 16512 3850 16522
rect 3976 16512 4042 16522
rect 4168 16512 4234 16522
rect 4360 16512 4426 16522
rect 4552 16512 4618 16522
rect 4744 16512 4810 16522
rect 4936 16512 5002 16522
rect 5128 16512 5184 16522
rect 5612 16512 5678 16522
rect 5804 16512 5870 16522
rect 5996 16512 6062 16522
rect 6188 16512 6254 16522
rect 6380 16512 6446 16522
rect 6572 16512 6638 16522
rect 6764 16512 6830 16522
rect 6956 16512 7012 16522
rect 7440 16512 7506 16522
rect 7632 16512 7698 16522
rect 7824 16512 7890 16522
rect 8016 16512 8082 16522
rect 8208 16512 8274 16522
rect 8400 16512 8466 16522
rect 8592 16512 8658 16522
rect 8784 16512 8840 16522
rect 9268 16512 9334 16522
rect 9460 16512 9526 16522
rect 9652 16512 9718 16522
rect 9844 16512 9910 16522
rect 10036 16512 10102 16522
rect 10228 16512 10294 16522
rect 10420 16512 10486 16522
rect 10612 16512 10668 16522
rect 11096 16512 11162 16522
rect 11288 16512 11354 16522
rect 11480 16512 11546 16522
rect 11672 16512 11738 16522
rect 11864 16512 11930 16522
rect 12056 16512 12122 16522
rect 12248 16512 12314 16522
rect 12440 16512 12496 16522
rect 12924 16512 12990 16522
rect 13116 16512 13182 16522
rect 13308 16512 13374 16522
rect 13500 16512 13566 16522
rect 13692 16512 13758 16522
rect 13884 16512 13950 16522
rect 14076 16512 14142 16522
rect 14268 16512 14324 16522
rect 14752 16512 14818 16522
rect 14944 16512 15010 16522
rect 15136 16512 15202 16522
rect 15328 16512 15394 16522
rect 15520 16512 15586 16522
rect 15712 16512 15778 16522
rect 15904 16512 15970 16522
rect 16096 16512 16152 16522
rect 16580 16512 16646 16522
rect 16772 16512 16838 16522
rect 16964 16512 17030 16522
rect 17156 16512 17222 16522
rect 17348 16512 17414 16522
rect 17540 16512 17606 16522
rect 17732 16512 17798 16522
rect 17924 16512 17980 16522
rect 18408 16512 18474 16522
rect 18600 16512 18666 16522
rect 18792 16512 18858 16522
rect 18984 16512 19050 16522
rect 19176 16512 19242 16522
rect 19368 16512 19434 16522
rect 19560 16512 19626 16522
rect 19752 16512 19808 16522
rect 20236 16512 20302 16522
rect 20428 16512 20494 16522
rect 20620 16512 20686 16522
rect 20812 16512 20878 16522
rect 21004 16512 21070 16522
rect 21196 16512 21262 16522
rect 21388 16512 21454 16522
rect 21580 16512 21636 16522
rect 32 16174 98 16184
rect 224 16174 290 16184
rect 416 16174 482 16184
rect 608 16174 674 16184
rect 800 16174 866 16184
rect 992 16174 1058 16184
rect 1184 16174 1250 16184
rect 1376 16174 1442 16184
rect 1860 16174 1926 16184
rect 2052 16174 2118 16184
rect 2244 16174 2310 16184
rect 2436 16174 2502 16184
rect 2628 16174 2694 16184
rect 2820 16174 2886 16184
rect 3012 16174 3078 16184
rect 3204 16174 3270 16184
rect 3688 16174 3754 16184
rect 3880 16174 3946 16184
rect 4072 16174 4138 16184
rect 4264 16174 4330 16184
rect 4456 16174 4522 16184
rect 4648 16174 4714 16184
rect 4840 16174 4906 16184
rect 5032 16174 5098 16184
rect 5516 16174 5582 16184
rect 5708 16174 5774 16184
rect 5900 16174 5966 16184
rect 6092 16174 6158 16184
rect 6284 16174 6350 16184
rect 6476 16174 6542 16184
rect 6668 16174 6734 16184
rect 6860 16174 6926 16184
rect 7344 16174 7410 16184
rect 7536 16174 7602 16184
rect 7728 16174 7794 16184
rect 7920 16174 7986 16184
rect 8112 16174 8178 16184
rect 8304 16174 8370 16184
rect 8496 16174 8562 16184
rect 8688 16174 8754 16184
rect 9172 16174 9238 16184
rect 9364 16174 9430 16184
rect 9556 16174 9622 16184
rect 9748 16174 9814 16184
rect 9940 16174 10006 16184
rect 10132 16174 10198 16184
rect 10324 16174 10390 16184
rect 10516 16174 10582 16184
rect 11000 16174 11066 16184
rect 11192 16174 11258 16184
rect 11384 16174 11450 16184
rect 11576 16174 11642 16184
rect 11768 16174 11834 16184
rect 11960 16174 12026 16184
rect 12152 16174 12218 16184
rect 12344 16174 12410 16184
rect 12828 16174 12894 16184
rect 13020 16174 13086 16184
rect 13212 16174 13278 16184
rect 13404 16174 13470 16184
rect 13596 16174 13662 16184
rect 13788 16174 13854 16184
rect 13980 16174 14046 16184
rect 14172 16174 14238 16184
rect 14656 16174 14722 16184
rect 14848 16174 14914 16184
rect 15040 16174 15106 16184
rect 15232 16174 15298 16184
rect 15424 16174 15490 16184
rect 15616 16174 15682 16184
rect 15808 16174 15874 16184
rect 16000 16174 16066 16184
rect 16484 16174 16550 16184
rect 16676 16174 16742 16184
rect 16868 16174 16934 16184
rect 17060 16174 17126 16184
rect 17252 16174 17318 16184
rect 17444 16174 17510 16184
rect 17636 16174 17702 16184
rect 17828 16174 17894 16184
rect 18312 16174 18378 16184
rect 18504 16174 18570 16184
rect 18696 16174 18762 16184
rect 18888 16174 18954 16184
rect 19080 16174 19146 16184
rect 19272 16174 19338 16184
rect 19464 16174 19530 16184
rect 19656 16174 19722 16184
rect 20140 16174 20206 16184
rect 20332 16174 20398 16184
rect 20524 16174 20590 16184
rect 20716 16174 20782 16184
rect 20908 16174 20974 16184
rect 21100 16174 21166 16184
rect 21292 16174 21358 16184
rect 21484 16174 21550 16184
rect 0 16021 32 16174
rect 98 16021 224 16174
rect 290 16021 416 16174
rect 482 16021 608 16174
rect 674 16021 800 16174
rect 866 16021 992 16174
rect 1058 16021 1184 16174
rect 1250 16021 1376 16174
rect 1828 16021 1860 16174
rect 1926 16021 2052 16174
rect 2118 16021 2244 16174
rect 2310 16021 2436 16174
rect 2502 16021 2628 16174
rect 2694 16021 2820 16174
rect 2886 16021 3012 16174
rect 3078 16021 3204 16174
rect 3656 16021 3688 16174
rect 3754 16021 3880 16174
rect 3946 16021 4072 16174
rect 4138 16021 4264 16174
rect 4330 16021 4456 16174
rect 4522 16021 4648 16174
rect 4714 16021 4840 16174
rect 4906 16021 5032 16174
rect 5484 16021 5516 16174
rect 5582 16021 5708 16174
rect 5774 16021 5900 16174
rect 5966 16021 6092 16174
rect 6158 16021 6284 16174
rect 6350 16021 6476 16174
rect 6542 16021 6668 16174
rect 6734 16021 6860 16174
rect 7312 16021 7344 16174
rect 7410 16021 7536 16174
rect 7602 16021 7728 16174
rect 7794 16021 7920 16174
rect 7986 16021 8112 16174
rect 8178 16021 8304 16174
rect 8370 16021 8496 16174
rect 8562 16021 8688 16174
rect 9140 16021 9172 16174
rect 9238 16021 9364 16174
rect 9430 16021 9556 16174
rect 9622 16021 9748 16174
rect 9814 16021 9940 16174
rect 10006 16021 10132 16174
rect 10198 16021 10324 16174
rect 10390 16021 10516 16174
rect 10968 16021 11000 16174
rect 11066 16021 11192 16174
rect 11258 16021 11384 16174
rect 11450 16021 11576 16174
rect 11642 16021 11768 16174
rect 11834 16021 11960 16174
rect 12026 16021 12152 16174
rect 12218 16021 12344 16174
rect 12796 16021 12828 16174
rect 12894 16021 13020 16174
rect 13086 16021 13212 16174
rect 13278 16021 13404 16174
rect 13470 16021 13596 16174
rect 13662 16021 13788 16174
rect 13854 16021 13980 16174
rect 14046 16021 14172 16174
rect 14624 16021 14656 16174
rect 14722 16021 14848 16174
rect 14914 16021 15040 16174
rect 15106 16021 15232 16174
rect 15298 16021 15424 16174
rect 15490 16021 15616 16174
rect 15682 16021 15808 16174
rect 15874 16021 16000 16174
rect 16452 16021 16484 16174
rect 16550 16021 16676 16174
rect 16742 16021 16868 16174
rect 16934 16021 17060 16174
rect 17126 16021 17252 16174
rect 17318 16021 17444 16174
rect 17510 16021 17636 16174
rect 17702 16021 17828 16174
rect 18280 16021 18312 16174
rect 18378 16021 18504 16174
rect 18570 16021 18696 16174
rect 18762 16021 18888 16174
rect 18954 16021 19080 16174
rect 19146 16021 19272 16174
rect 19338 16021 19464 16174
rect 19530 16021 19656 16174
rect 20108 16021 20140 16174
rect 20206 16021 20332 16174
rect 20398 16021 20524 16174
rect 20590 16021 20716 16174
rect 20782 16021 20908 16174
rect 20974 16021 21100 16174
rect 21166 16021 21292 16174
rect 21358 16021 21484 16174
rect 32 16011 98 16021
rect 224 16011 290 16021
rect 416 16011 482 16021
rect 608 16011 674 16021
rect 800 16011 866 16021
rect 992 16011 1058 16021
rect 1184 16011 1250 16021
rect 1376 16011 1442 16021
rect 1860 16011 1926 16021
rect 2052 16011 2118 16021
rect 2244 16011 2310 16021
rect 2436 16011 2502 16021
rect 2628 16011 2694 16021
rect 2820 16011 2886 16021
rect 3012 16011 3078 16021
rect 3204 16011 3270 16021
rect 3688 16011 3754 16021
rect 3880 16011 3946 16021
rect 4072 16011 4138 16021
rect 4264 16011 4330 16021
rect 4456 16011 4522 16021
rect 4648 16011 4714 16021
rect 4840 16011 4906 16021
rect 5032 16011 5098 16021
rect 5516 16011 5582 16021
rect 5708 16011 5774 16021
rect 5900 16011 5966 16021
rect 6092 16011 6158 16021
rect 6284 16011 6350 16021
rect 6476 16011 6542 16021
rect 6668 16011 6734 16021
rect 6860 16011 6926 16021
rect 7344 16011 7410 16021
rect 7536 16011 7602 16021
rect 7728 16011 7794 16021
rect 7920 16011 7986 16021
rect 8112 16011 8178 16021
rect 8304 16011 8370 16021
rect 8496 16011 8562 16021
rect 8688 16011 8754 16021
rect 9172 16011 9238 16021
rect 9364 16011 9430 16021
rect 9556 16011 9622 16021
rect 9748 16011 9814 16021
rect 9940 16011 10006 16021
rect 10132 16011 10198 16021
rect 10324 16011 10390 16021
rect 10516 16011 10582 16021
rect 11000 16011 11066 16021
rect 11192 16011 11258 16021
rect 11384 16011 11450 16021
rect 11576 16011 11642 16021
rect 11768 16011 11834 16021
rect 11960 16011 12026 16021
rect 12152 16011 12218 16021
rect 12344 16011 12410 16021
rect 12828 16011 12894 16021
rect 13020 16011 13086 16021
rect 13212 16011 13278 16021
rect 13404 16011 13470 16021
rect 13596 16011 13662 16021
rect 13788 16011 13854 16021
rect 13980 16011 14046 16021
rect 14172 16011 14238 16021
rect 14656 16011 14722 16021
rect 14848 16011 14914 16021
rect 15040 16011 15106 16021
rect 15232 16011 15298 16021
rect 15424 16011 15490 16021
rect 15616 16011 15682 16021
rect 15808 16011 15874 16021
rect 16000 16011 16066 16021
rect 16484 16011 16550 16021
rect 16676 16011 16742 16021
rect 16868 16011 16934 16021
rect 17060 16011 17126 16021
rect 17252 16011 17318 16021
rect 17444 16011 17510 16021
rect 17636 16011 17702 16021
rect 17828 16011 17894 16021
rect 18312 16011 18378 16021
rect 18504 16011 18570 16021
rect 18696 16011 18762 16021
rect 18888 16011 18954 16021
rect 19080 16011 19146 16021
rect 19272 16011 19338 16021
rect 19464 16011 19530 16021
rect 19656 16011 19722 16021
rect 20140 16011 20206 16021
rect 20332 16011 20398 16021
rect 20524 16011 20590 16021
rect 20716 16011 20782 16021
rect 20908 16011 20974 16021
rect 21100 16011 21166 16021
rect 21292 16011 21358 16021
rect 21484 16011 21550 16021
rect 128 15961 194 15971
rect 320 15961 386 15971
rect 512 15961 578 15971
rect 704 15961 770 15971
rect 896 15961 962 15971
rect 1088 15961 1154 15971
rect 1280 15961 1346 15971
rect 1472 15961 1528 15971
rect 1956 15961 2022 15971
rect 2148 15961 2214 15971
rect 2340 15961 2406 15971
rect 2532 15961 2598 15971
rect 2724 15961 2790 15971
rect 2916 15961 2982 15971
rect 3108 15961 3174 15971
rect 3300 15961 3356 15971
rect 3784 15961 3850 15971
rect 3976 15961 4042 15971
rect 4168 15961 4234 15971
rect 4360 15961 4426 15971
rect 4552 15961 4618 15971
rect 4744 15961 4810 15971
rect 4936 15961 5002 15971
rect 5128 15961 5184 15971
rect 5612 15961 5678 15971
rect 5804 15961 5870 15971
rect 5996 15961 6062 15971
rect 6188 15961 6254 15971
rect 6380 15961 6446 15971
rect 6572 15961 6638 15971
rect 6764 15961 6830 15971
rect 6956 15961 7012 15971
rect 7440 15961 7506 15971
rect 7632 15961 7698 15971
rect 7824 15961 7890 15971
rect 8016 15961 8082 15971
rect 8208 15961 8274 15971
rect 8400 15961 8466 15971
rect 8592 15961 8658 15971
rect 8784 15961 8840 15971
rect 9268 15961 9334 15971
rect 9460 15961 9526 15971
rect 9652 15961 9718 15971
rect 9844 15961 9910 15971
rect 10036 15961 10102 15971
rect 10228 15961 10294 15971
rect 10420 15961 10486 15971
rect 10612 15961 10668 15971
rect 11096 15961 11162 15971
rect 11288 15961 11354 15971
rect 11480 15961 11546 15971
rect 11672 15961 11738 15971
rect 11864 15961 11930 15971
rect 12056 15961 12122 15971
rect 12248 15961 12314 15971
rect 12440 15961 12496 15971
rect 12924 15961 12990 15971
rect 13116 15961 13182 15971
rect 13308 15961 13374 15971
rect 13500 15961 13566 15971
rect 13692 15961 13758 15971
rect 13884 15961 13950 15971
rect 14076 15961 14142 15971
rect 14268 15961 14324 15971
rect 14752 15961 14818 15971
rect 14944 15961 15010 15971
rect 15136 15961 15202 15971
rect 15328 15961 15394 15971
rect 15520 15961 15586 15971
rect 15712 15961 15778 15971
rect 15904 15961 15970 15971
rect 16096 15961 16152 15971
rect 16580 15961 16646 15971
rect 16772 15961 16838 15971
rect 16964 15961 17030 15971
rect 17156 15961 17222 15971
rect 17348 15961 17414 15971
rect 17540 15961 17606 15971
rect 17732 15961 17798 15971
rect 17924 15961 17980 15971
rect 18408 15961 18474 15971
rect 18600 15961 18666 15971
rect 18792 15961 18858 15971
rect 18984 15961 19050 15971
rect 19176 15961 19242 15971
rect 19368 15961 19434 15971
rect 19560 15961 19626 15971
rect 19752 15961 19808 15971
rect 20236 15961 20302 15971
rect 20428 15961 20494 15971
rect 20620 15961 20686 15971
rect 20812 15961 20878 15971
rect 21004 15961 21070 15971
rect 21196 15961 21262 15971
rect 21388 15961 21454 15971
rect 21580 15961 21636 15971
rect 0 15808 128 15961
rect 194 15808 320 15961
rect 386 15808 512 15961
rect 578 15808 704 15961
rect 770 15808 896 15961
rect 962 15808 1088 15961
rect 1154 15808 1280 15961
rect 1346 15808 1472 15961
rect 1528 15808 1708 15961
rect 1828 15808 1956 15961
rect 2022 15808 2148 15961
rect 2214 15808 2340 15961
rect 2406 15808 2532 15961
rect 2598 15808 2724 15961
rect 2790 15808 2916 15961
rect 2982 15808 3108 15961
rect 3174 15808 3300 15961
rect 3356 15808 3536 15961
rect 3656 15808 3784 15961
rect 3850 15808 3976 15961
rect 4042 15808 4168 15961
rect 4234 15808 4360 15961
rect 4426 15808 4552 15961
rect 4618 15808 4744 15961
rect 4810 15808 4936 15961
rect 5002 15808 5128 15961
rect 5184 15808 5364 15961
rect 5484 15808 5612 15961
rect 5678 15808 5804 15961
rect 5870 15808 5996 15961
rect 6062 15808 6188 15961
rect 6254 15808 6380 15961
rect 6446 15808 6572 15961
rect 6638 15808 6764 15961
rect 6830 15808 6956 15961
rect 7012 15808 7192 15961
rect 7312 15808 7440 15961
rect 7506 15808 7632 15961
rect 7698 15808 7824 15961
rect 7890 15808 8016 15961
rect 8082 15808 8208 15961
rect 8274 15808 8400 15961
rect 8466 15808 8592 15961
rect 8658 15808 8784 15961
rect 8840 15808 9020 15961
rect 9140 15808 9268 15961
rect 9334 15808 9460 15961
rect 9526 15808 9652 15961
rect 9718 15808 9844 15961
rect 9910 15808 10036 15961
rect 10102 15808 10228 15961
rect 10294 15808 10420 15961
rect 10486 15808 10612 15961
rect 10668 15808 10848 15961
rect 10968 15808 11096 15961
rect 11162 15808 11288 15961
rect 11354 15808 11480 15961
rect 11546 15808 11672 15961
rect 11738 15808 11864 15961
rect 11930 15808 12056 15961
rect 12122 15808 12248 15961
rect 12314 15808 12440 15961
rect 12496 15808 12676 15961
rect 12796 15808 12924 15961
rect 12990 15808 13116 15961
rect 13182 15808 13308 15961
rect 13374 15808 13500 15961
rect 13566 15808 13692 15961
rect 13758 15808 13884 15961
rect 13950 15808 14076 15961
rect 14142 15808 14268 15961
rect 14324 15808 14504 15961
rect 14624 15808 14752 15961
rect 14818 15808 14944 15961
rect 15010 15808 15136 15961
rect 15202 15808 15328 15961
rect 15394 15808 15520 15961
rect 15586 15808 15712 15961
rect 15778 15808 15904 15961
rect 15970 15808 16096 15961
rect 16152 15808 16332 15961
rect 16452 15808 16580 15961
rect 16646 15808 16772 15961
rect 16838 15808 16964 15961
rect 17030 15808 17156 15961
rect 17222 15808 17348 15961
rect 17414 15808 17540 15961
rect 17606 15808 17732 15961
rect 17798 15808 17924 15961
rect 17980 15808 18160 15961
rect 18280 15808 18408 15961
rect 18474 15808 18600 15961
rect 18666 15808 18792 15961
rect 18858 15808 18984 15961
rect 19050 15808 19176 15961
rect 19242 15808 19368 15961
rect 19434 15808 19560 15961
rect 19626 15808 19752 15961
rect 19808 15808 19988 15961
rect 20108 15808 20236 15961
rect 20302 15808 20428 15961
rect 20494 15808 20620 15961
rect 20686 15808 20812 15961
rect 20878 15808 21004 15961
rect 21070 15808 21196 15961
rect 21262 15808 21388 15961
rect 21454 15808 21580 15961
rect 21636 15808 21816 15961
rect 128 15798 194 15808
rect 320 15798 386 15808
rect 512 15798 578 15808
rect 704 15798 770 15808
rect 896 15798 962 15808
rect 1088 15798 1154 15808
rect 1280 15798 1346 15808
rect 1472 15798 1528 15808
rect 1956 15798 2022 15808
rect 2148 15798 2214 15808
rect 2340 15798 2406 15808
rect 2532 15798 2598 15808
rect 2724 15798 2790 15808
rect 2916 15798 2982 15808
rect 3108 15798 3174 15808
rect 3300 15798 3356 15808
rect 3784 15798 3850 15808
rect 3976 15798 4042 15808
rect 4168 15798 4234 15808
rect 4360 15798 4426 15808
rect 4552 15798 4618 15808
rect 4744 15798 4810 15808
rect 4936 15798 5002 15808
rect 5128 15798 5184 15808
rect 5612 15798 5678 15808
rect 5804 15798 5870 15808
rect 5996 15798 6062 15808
rect 6188 15798 6254 15808
rect 6380 15798 6446 15808
rect 6572 15798 6638 15808
rect 6764 15798 6830 15808
rect 6956 15798 7012 15808
rect 7440 15798 7506 15808
rect 7632 15798 7698 15808
rect 7824 15798 7890 15808
rect 8016 15798 8082 15808
rect 8208 15798 8274 15808
rect 8400 15798 8466 15808
rect 8592 15798 8658 15808
rect 8784 15798 8840 15808
rect 9268 15798 9334 15808
rect 9460 15798 9526 15808
rect 9652 15798 9718 15808
rect 9844 15798 9910 15808
rect 10036 15798 10102 15808
rect 10228 15798 10294 15808
rect 10420 15798 10486 15808
rect 10612 15798 10668 15808
rect 11096 15798 11162 15808
rect 11288 15798 11354 15808
rect 11480 15798 11546 15808
rect 11672 15798 11738 15808
rect 11864 15798 11930 15808
rect 12056 15798 12122 15808
rect 12248 15798 12314 15808
rect 12440 15798 12496 15808
rect 12924 15798 12990 15808
rect 13116 15798 13182 15808
rect 13308 15798 13374 15808
rect 13500 15798 13566 15808
rect 13692 15798 13758 15808
rect 13884 15798 13950 15808
rect 14076 15798 14142 15808
rect 14268 15798 14324 15808
rect 14752 15798 14818 15808
rect 14944 15798 15010 15808
rect 15136 15798 15202 15808
rect 15328 15798 15394 15808
rect 15520 15798 15586 15808
rect 15712 15798 15778 15808
rect 15904 15798 15970 15808
rect 16096 15798 16152 15808
rect 16580 15798 16646 15808
rect 16772 15798 16838 15808
rect 16964 15798 17030 15808
rect 17156 15798 17222 15808
rect 17348 15798 17414 15808
rect 17540 15798 17606 15808
rect 17732 15798 17798 15808
rect 17924 15798 17980 15808
rect 18408 15798 18474 15808
rect 18600 15798 18666 15808
rect 18792 15798 18858 15808
rect 18984 15798 19050 15808
rect 19176 15798 19242 15808
rect 19368 15798 19434 15808
rect 19560 15798 19626 15808
rect 19752 15798 19808 15808
rect 20236 15798 20302 15808
rect 20428 15798 20494 15808
rect 20620 15798 20686 15808
rect 20812 15798 20878 15808
rect 21004 15798 21070 15808
rect 21196 15798 21262 15808
rect 21388 15798 21454 15808
rect 21580 15798 21636 15808
rect 32 15460 98 15470
rect 224 15460 290 15470
rect 416 15460 482 15470
rect 608 15460 674 15470
rect 800 15460 866 15470
rect 992 15460 1058 15470
rect 1184 15460 1250 15470
rect 1376 15460 1442 15470
rect 1860 15460 1926 15470
rect 2052 15460 2118 15470
rect 2244 15460 2310 15470
rect 2436 15460 2502 15470
rect 2628 15460 2694 15470
rect 2820 15460 2886 15470
rect 3012 15460 3078 15470
rect 3204 15460 3270 15470
rect 3688 15460 3754 15470
rect 3880 15460 3946 15470
rect 4072 15460 4138 15470
rect 4264 15460 4330 15470
rect 4456 15460 4522 15470
rect 4648 15460 4714 15470
rect 4840 15460 4906 15470
rect 5032 15460 5098 15470
rect 5516 15460 5582 15470
rect 5708 15460 5774 15470
rect 5900 15460 5966 15470
rect 6092 15460 6158 15470
rect 6284 15460 6350 15470
rect 6476 15460 6542 15470
rect 6668 15460 6734 15470
rect 6860 15460 6926 15470
rect 7344 15460 7410 15470
rect 7536 15460 7602 15470
rect 7728 15460 7794 15470
rect 7920 15460 7986 15470
rect 8112 15460 8178 15470
rect 8304 15460 8370 15470
rect 8496 15460 8562 15470
rect 8688 15460 8754 15470
rect 9172 15460 9238 15470
rect 9364 15460 9430 15470
rect 9556 15460 9622 15470
rect 9748 15460 9814 15470
rect 9940 15460 10006 15470
rect 10132 15460 10198 15470
rect 10324 15460 10390 15470
rect 10516 15460 10582 15470
rect 11000 15460 11066 15470
rect 11192 15460 11258 15470
rect 11384 15460 11450 15470
rect 11576 15460 11642 15470
rect 11768 15460 11834 15470
rect 11960 15460 12026 15470
rect 12152 15460 12218 15470
rect 12344 15460 12410 15470
rect 12828 15460 12894 15470
rect 13020 15460 13086 15470
rect 13212 15460 13278 15470
rect 13404 15460 13470 15470
rect 13596 15460 13662 15470
rect 13788 15460 13854 15470
rect 13980 15460 14046 15470
rect 14172 15460 14238 15470
rect 14656 15460 14722 15470
rect 14848 15460 14914 15470
rect 15040 15460 15106 15470
rect 15232 15460 15298 15470
rect 15424 15460 15490 15470
rect 15616 15460 15682 15470
rect 15808 15460 15874 15470
rect 16000 15460 16066 15470
rect 16484 15460 16550 15470
rect 16676 15460 16742 15470
rect 16868 15460 16934 15470
rect 17060 15460 17126 15470
rect 17252 15460 17318 15470
rect 17444 15460 17510 15470
rect 17636 15460 17702 15470
rect 17828 15460 17894 15470
rect 18312 15460 18378 15470
rect 18504 15460 18570 15470
rect 18696 15460 18762 15470
rect 18888 15460 18954 15470
rect 19080 15460 19146 15470
rect 19272 15460 19338 15470
rect 19464 15460 19530 15470
rect 19656 15460 19722 15470
rect 20140 15460 20206 15470
rect 20332 15460 20398 15470
rect 20524 15460 20590 15470
rect 20716 15460 20782 15470
rect 20908 15460 20974 15470
rect 21100 15460 21166 15470
rect 21292 15460 21358 15470
rect 21484 15460 21550 15470
rect 0 15307 32 15460
rect 98 15307 224 15460
rect 290 15307 416 15460
rect 482 15307 608 15460
rect 674 15307 800 15460
rect 866 15307 992 15460
rect 1058 15307 1184 15460
rect 1250 15307 1376 15460
rect 1828 15307 1860 15460
rect 1926 15307 2052 15460
rect 2118 15307 2244 15460
rect 2310 15307 2436 15460
rect 2502 15307 2628 15460
rect 2694 15307 2820 15460
rect 2886 15307 3012 15460
rect 3078 15307 3204 15460
rect 3656 15307 3688 15460
rect 3754 15307 3880 15460
rect 3946 15307 4072 15460
rect 4138 15307 4264 15460
rect 4330 15307 4456 15460
rect 4522 15307 4648 15460
rect 4714 15307 4840 15460
rect 4906 15307 5032 15460
rect 5484 15307 5516 15460
rect 5582 15307 5708 15460
rect 5774 15307 5900 15460
rect 5966 15307 6092 15460
rect 6158 15307 6284 15460
rect 6350 15307 6476 15460
rect 6542 15307 6668 15460
rect 6734 15307 6860 15460
rect 7312 15307 7344 15460
rect 7410 15307 7536 15460
rect 7602 15307 7728 15460
rect 7794 15307 7920 15460
rect 7986 15307 8112 15460
rect 8178 15307 8304 15460
rect 8370 15307 8496 15460
rect 8562 15307 8688 15460
rect 9140 15307 9172 15460
rect 9238 15307 9364 15460
rect 9430 15307 9556 15460
rect 9622 15307 9748 15460
rect 9814 15307 9940 15460
rect 10006 15307 10132 15460
rect 10198 15307 10324 15460
rect 10390 15307 10516 15460
rect 10968 15307 11000 15460
rect 11066 15307 11192 15460
rect 11258 15307 11384 15460
rect 11450 15307 11576 15460
rect 11642 15307 11768 15460
rect 11834 15307 11960 15460
rect 12026 15307 12152 15460
rect 12218 15307 12344 15460
rect 12796 15307 12828 15460
rect 12894 15307 13020 15460
rect 13086 15307 13212 15460
rect 13278 15307 13404 15460
rect 13470 15307 13596 15460
rect 13662 15307 13788 15460
rect 13854 15307 13980 15460
rect 14046 15307 14172 15460
rect 14624 15307 14656 15460
rect 14722 15307 14848 15460
rect 14914 15307 15040 15460
rect 15106 15307 15232 15460
rect 15298 15307 15424 15460
rect 15490 15307 15616 15460
rect 15682 15307 15808 15460
rect 15874 15307 16000 15460
rect 16452 15307 16484 15460
rect 16550 15307 16676 15460
rect 16742 15307 16868 15460
rect 16934 15307 17060 15460
rect 17126 15307 17252 15460
rect 17318 15307 17444 15460
rect 17510 15307 17636 15460
rect 17702 15307 17828 15460
rect 18280 15307 18312 15460
rect 18378 15307 18504 15460
rect 18570 15307 18696 15460
rect 18762 15307 18888 15460
rect 18954 15307 19080 15460
rect 19146 15307 19272 15460
rect 19338 15307 19464 15460
rect 19530 15307 19656 15460
rect 20108 15307 20140 15460
rect 20206 15307 20332 15460
rect 20398 15307 20524 15460
rect 20590 15307 20716 15460
rect 20782 15307 20908 15460
rect 20974 15307 21100 15460
rect 21166 15307 21292 15460
rect 21358 15307 21484 15460
rect 32 15297 98 15307
rect 224 15297 290 15307
rect 416 15297 482 15307
rect 608 15297 674 15307
rect 800 15297 866 15307
rect 992 15297 1058 15307
rect 1184 15297 1250 15307
rect 1376 15297 1442 15307
rect 1860 15297 1926 15307
rect 2052 15297 2118 15307
rect 2244 15297 2310 15307
rect 2436 15297 2502 15307
rect 2628 15297 2694 15307
rect 2820 15297 2886 15307
rect 3012 15297 3078 15307
rect 3204 15297 3270 15307
rect 3688 15297 3754 15307
rect 3880 15297 3946 15307
rect 4072 15297 4138 15307
rect 4264 15297 4330 15307
rect 4456 15297 4522 15307
rect 4648 15297 4714 15307
rect 4840 15297 4906 15307
rect 5032 15297 5098 15307
rect 5516 15297 5582 15307
rect 5708 15297 5774 15307
rect 5900 15297 5966 15307
rect 6092 15297 6158 15307
rect 6284 15297 6350 15307
rect 6476 15297 6542 15307
rect 6668 15297 6734 15307
rect 6860 15297 6926 15307
rect 7344 15297 7410 15307
rect 7536 15297 7602 15307
rect 7728 15297 7794 15307
rect 7920 15297 7986 15307
rect 8112 15297 8178 15307
rect 8304 15297 8370 15307
rect 8496 15297 8562 15307
rect 8688 15297 8754 15307
rect 9172 15297 9238 15307
rect 9364 15297 9430 15307
rect 9556 15297 9622 15307
rect 9748 15297 9814 15307
rect 9940 15297 10006 15307
rect 10132 15297 10198 15307
rect 10324 15297 10390 15307
rect 10516 15297 10582 15307
rect 11000 15297 11066 15307
rect 11192 15297 11258 15307
rect 11384 15297 11450 15307
rect 11576 15297 11642 15307
rect 11768 15297 11834 15307
rect 11960 15297 12026 15307
rect 12152 15297 12218 15307
rect 12344 15297 12410 15307
rect 12828 15297 12894 15307
rect 13020 15297 13086 15307
rect 13212 15297 13278 15307
rect 13404 15297 13470 15307
rect 13596 15297 13662 15307
rect 13788 15297 13854 15307
rect 13980 15297 14046 15307
rect 14172 15297 14238 15307
rect 14656 15297 14722 15307
rect 14848 15297 14914 15307
rect 15040 15297 15106 15307
rect 15232 15297 15298 15307
rect 15424 15297 15490 15307
rect 15616 15297 15682 15307
rect 15808 15297 15874 15307
rect 16000 15297 16066 15307
rect 16484 15297 16550 15307
rect 16676 15297 16742 15307
rect 16868 15297 16934 15307
rect 17060 15297 17126 15307
rect 17252 15297 17318 15307
rect 17444 15297 17510 15307
rect 17636 15297 17702 15307
rect 17828 15297 17894 15307
rect 18312 15297 18378 15307
rect 18504 15297 18570 15307
rect 18696 15297 18762 15307
rect 18888 15297 18954 15307
rect 19080 15297 19146 15307
rect 19272 15297 19338 15307
rect 19464 15297 19530 15307
rect 19656 15297 19722 15307
rect 20140 15297 20206 15307
rect 20332 15297 20398 15307
rect 20524 15297 20590 15307
rect 20716 15297 20782 15307
rect 20908 15297 20974 15307
rect 21100 15297 21166 15307
rect 21292 15297 21358 15307
rect 21484 15297 21550 15307
rect 128 15247 194 15257
rect 320 15247 386 15257
rect 512 15247 578 15257
rect 704 15247 770 15257
rect 896 15247 962 15257
rect 1088 15247 1154 15257
rect 1280 15247 1346 15257
rect 1472 15247 1528 15257
rect 1956 15247 2022 15257
rect 2148 15247 2214 15257
rect 2340 15247 2406 15257
rect 2532 15247 2598 15257
rect 2724 15247 2790 15257
rect 2916 15247 2982 15257
rect 3108 15247 3174 15257
rect 3300 15247 3356 15257
rect 3784 15247 3850 15257
rect 3976 15247 4042 15257
rect 4168 15247 4234 15257
rect 4360 15247 4426 15257
rect 4552 15247 4618 15257
rect 4744 15247 4810 15257
rect 4936 15247 5002 15257
rect 5128 15247 5184 15257
rect 5612 15247 5678 15257
rect 5804 15247 5870 15257
rect 5996 15247 6062 15257
rect 6188 15247 6254 15257
rect 6380 15247 6446 15257
rect 6572 15247 6638 15257
rect 6764 15247 6830 15257
rect 6956 15247 7012 15257
rect 7440 15247 7506 15257
rect 7632 15247 7698 15257
rect 7824 15247 7890 15257
rect 8016 15247 8082 15257
rect 8208 15247 8274 15257
rect 8400 15247 8466 15257
rect 8592 15247 8658 15257
rect 8784 15247 8840 15257
rect 9268 15247 9334 15257
rect 9460 15247 9526 15257
rect 9652 15247 9718 15257
rect 9844 15247 9910 15257
rect 10036 15247 10102 15257
rect 10228 15247 10294 15257
rect 10420 15247 10486 15257
rect 10612 15247 10668 15257
rect 11096 15247 11162 15257
rect 11288 15247 11354 15257
rect 11480 15247 11546 15257
rect 11672 15247 11738 15257
rect 11864 15247 11930 15257
rect 12056 15247 12122 15257
rect 12248 15247 12314 15257
rect 12440 15247 12496 15257
rect 12924 15247 12990 15257
rect 13116 15247 13182 15257
rect 13308 15247 13374 15257
rect 13500 15247 13566 15257
rect 13692 15247 13758 15257
rect 13884 15247 13950 15257
rect 14076 15247 14142 15257
rect 14268 15247 14324 15257
rect 14752 15247 14818 15257
rect 14944 15247 15010 15257
rect 15136 15247 15202 15257
rect 15328 15247 15394 15257
rect 15520 15247 15586 15257
rect 15712 15247 15778 15257
rect 15904 15247 15970 15257
rect 16096 15247 16152 15257
rect 16580 15247 16646 15257
rect 16772 15247 16838 15257
rect 16964 15247 17030 15257
rect 17156 15247 17222 15257
rect 17348 15247 17414 15257
rect 17540 15247 17606 15257
rect 17732 15247 17798 15257
rect 17924 15247 17980 15257
rect 18408 15247 18474 15257
rect 18600 15247 18666 15257
rect 18792 15247 18858 15257
rect 18984 15247 19050 15257
rect 19176 15247 19242 15257
rect 19368 15247 19434 15257
rect 19560 15247 19626 15257
rect 19752 15247 19808 15257
rect 20236 15247 20302 15257
rect 20428 15247 20494 15257
rect 20620 15247 20686 15257
rect 20812 15247 20878 15257
rect 21004 15247 21070 15257
rect 21196 15247 21262 15257
rect 21388 15247 21454 15257
rect 21580 15247 21636 15257
rect 0 15094 128 15247
rect 194 15094 320 15247
rect 386 15094 512 15247
rect 578 15094 704 15247
rect 770 15094 896 15247
rect 962 15094 1088 15247
rect 1154 15094 1280 15247
rect 1346 15094 1472 15247
rect 1528 15094 1708 15247
rect 1828 15094 1956 15247
rect 2022 15094 2148 15247
rect 2214 15094 2340 15247
rect 2406 15094 2532 15247
rect 2598 15094 2724 15247
rect 2790 15094 2916 15247
rect 2982 15094 3108 15247
rect 3174 15094 3300 15247
rect 3356 15094 3536 15247
rect 3656 15094 3784 15247
rect 3850 15094 3976 15247
rect 4042 15094 4168 15247
rect 4234 15094 4360 15247
rect 4426 15094 4552 15247
rect 4618 15094 4744 15247
rect 4810 15094 4936 15247
rect 5002 15094 5128 15247
rect 5184 15094 5364 15247
rect 5484 15094 5612 15247
rect 5678 15094 5804 15247
rect 5870 15094 5996 15247
rect 6062 15094 6188 15247
rect 6254 15094 6380 15247
rect 6446 15094 6572 15247
rect 6638 15094 6764 15247
rect 6830 15094 6956 15247
rect 7012 15094 7192 15247
rect 7312 15094 7440 15247
rect 7506 15094 7632 15247
rect 7698 15094 7824 15247
rect 7890 15094 8016 15247
rect 8082 15094 8208 15247
rect 8274 15094 8400 15247
rect 8466 15094 8592 15247
rect 8658 15094 8784 15247
rect 8840 15094 9020 15247
rect 9140 15094 9268 15247
rect 9334 15094 9460 15247
rect 9526 15094 9652 15247
rect 9718 15094 9844 15247
rect 9910 15094 10036 15247
rect 10102 15094 10228 15247
rect 10294 15094 10420 15247
rect 10486 15094 10612 15247
rect 10668 15094 10848 15247
rect 10968 15094 11096 15247
rect 11162 15094 11288 15247
rect 11354 15094 11480 15247
rect 11546 15094 11672 15247
rect 11738 15094 11864 15247
rect 11930 15094 12056 15247
rect 12122 15094 12248 15247
rect 12314 15094 12440 15247
rect 12496 15094 12676 15247
rect 12796 15094 12924 15247
rect 12990 15094 13116 15247
rect 13182 15094 13308 15247
rect 13374 15094 13500 15247
rect 13566 15094 13692 15247
rect 13758 15094 13884 15247
rect 13950 15094 14076 15247
rect 14142 15094 14268 15247
rect 14324 15094 14504 15247
rect 14624 15094 14752 15247
rect 14818 15094 14944 15247
rect 15010 15094 15136 15247
rect 15202 15094 15328 15247
rect 15394 15094 15520 15247
rect 15586 15094 15712 15247
rect 15778 15094 15904 15247
rect 15970 15094 16096 15247
rect 16152 15094 16332 15247
rect 16452 15094 16580 15247
rect 16646 15094 16772 15247
rect 16838 15094 16964 15247
rect 17030 15094 17156 15247
rect 17222 15094 17348 15247
rect 17414 15094 17540 15247
rect 17606 15094 17732 15247
rect 17798 15094 17924 15247
rect 17980 15094 18160 15247
rect 18280 15094 18408 15247
rect 18474 15094 18600 15247
rect 18666 15094 18792 15247
rect 18858 15094 18984 15247
rect 19050 15094 19176 15247
rect 19242 15094 19368 15247
rect 19434 15094 19560 15247
rect 19626 15094 19752 15247
rect 19808 15094 19988 15247
rect 20108 15094 20236 15247
rect 20302 15094 20428 15247
rect 20494 15094 20620 15247
rect 20686 15094 20812 15247
rect 20878 15094 21004 15247
rect 21070 15094 21196 15247
rect 21262 15094 21388 15247
rect 21454 15094 21580 15247
rect 21636 15094 21816 15247
rect 128 15084 194 15094
rect 320 15084 386 15094
rect 512 15084 578 15094
rect 704 15084 770 15094
rect 896 15084 962 15094
rect 1088 15084 1154 15094
rect 1280 15084 1346 15094
rect 1472 15084 1528 15094
rect 1956 15084 2022 15094
rect 2148 15084 2214 15094
rect 2340 15084 2406 15094
rect 2532 15084 2598 15094
rect 2724 15084 2790 15094
rect 2916 15084 2982 15094
rect 3108 15084 3174 15094
rect 3300 15084 3356 15094
rect 3784 15084 3850 15094
rect 3976 15084 4042 15094
rect 4168 15084 4234 15094
rect 4360 15084 4426 15094
rect 4552 15084 4618 15094
rect 4744 15084 4810 15094
rect 4936 15084 5002 15094
rect 5128 15084 5184 15094
rect 5612 15084 5678 15094
rect 5804 15084 5870 15094
rect 5996 15084 6062 15094
rect 6188 15084 6254 15094
rect 6380 15084 6446 15094
rect 6572 15084 6638 15094
rect 6764 15084 6830 15094
rect 6956 15084 7012 15094
rect 7440 15084 7506 15094
rect 7632 15084 7698 15094
rect 7824 15084 7890 15094
rect 8016 15084 8082 15094
rect 8208 15084 8274 15094
rect 8400 15084 8466 15094
rect 8592 15084 8658 15094
rect 8784 15084 8840 15094
rect 9268 15084 9334 15094
rect 9460 15084 9526 15094
rect 9652 15084 9718 15094
rect 9844 15084 9910 15094
rect 10036 15084 10102 15094
rect 10228 15084 10294 15094
rect 10420 15084 10486 15094
rect 10612 15084 10668 15094
rect 11096 15084 11162 15094
rect 11288 15084 11354 15094
rect 11480 15084 11546 15094
rect 11672 15084 11738 15094
rect 11864 15084 11930 15094
rect 12056 15084 12122 15094
rect 12248 15084 12314 15094
rect 12440 15084 12496 15094
rect 12924 15084 12990 15094
rect 13116 15084 13182 15094
rect 13308 15084 13374 15094
rect 13500 15084 13566 15094
rect 13692 15084 13758 15094
rect 13884 15084 13950 15094
rect 14076 15084 14142 15094
rect 14268 15084 14324 15094
rect 14752 15084 14818 15094
rect 14944 15084 15010 15094
rect 15136 15084 15202 15094
rect 15328 15084 15394 15094
rect 15520 15084 15586 15094
rect 15712 15084 15778 15094
rect 15904 15084 15970 15094
rect 16096 15084 16152 15094
rect 16580 15084 16646 15094
rect 16772 15084 16838 15094
rect 16964 15084 17030 15094
rect 17156 15084 17222 15094
rect 17348 15084 17414 15094
rect 17540 15084 17606 15094
rect 17732 15084 17798 15094
rect 17924 15084 17980 15094
rect 18408 15084 18474 15094
rect 18600 15084 18666 15094
rect 18792 15084 18858 15094
rect 18984 15084 19050 15094
rect 19176 15084 19242 15094
rect 19368 15084 19434 15094
rect 19560 15084 19626 15094
rect 19752 15084 19808 15094
rect 20236 15084 20302 15094
rect 20428 15084 20494 15094
rect 20620 15084 20686 15094
rect 20812 15084 20878 15094
rect 21004 15084 21070 15094
rect 21196 15084 21262 15094
rect 21388 15084 21454 15094
rect 21580 15084 21636 15094
rect 32 14746 98 14756
rect 224 14746 290 14756
rect 416 14746 482 14756
rect 608 14746 674 14756
rect 800 14746 866 14756
rect 992 14746 1058 14756
rect 1184 14746 1250 14756
rect 1376 14746 1442 14756
rect 1860 14746 1926 14756
rect 2052 14746 2118 14756
rect 2244 14746 2310 14756
rect 2436 14746 2502 14756
rect 2628 14746 2694 14756
rect 2820 14746 2886 14756
rect 3012 14746 3078 14756
rect 3204 14746 3270 14756
rect 3688 14746 3754 14756
rect 3880 14746 3946 14756
rect 4072 14746 4138 14756
rect 4264 14746 4330 14756
rect 4456 14746 4522 14756
rect 4648 14746 4714 14756
rect 4840 14746 4906 14756
rect 5032 14746 5098 14756
rect 5516 14746 5582 14756
rect 5708 14746 5774 14756
rect 5900 14746 5966 14756
rect 6092 14746 6158 14756
rect 6284 14746 6350 14756
rect 6476 14746 6542 14756
rect 6668 14746 6734 14756
rect 6860 14746 6926 14756
rect 7344 14746 7410 14756
rect 7536 14746 7602 14756
rect 7728 14746 7794 14756
rect 7920 14746 7986 14756
rect 8112 14746 8178 14756
rect 8304 14746 8370 14756
rect 8496 14746 8562 14756
rect 8688 14746 8754 14756
rect 9172 14746 9238 14756
rect 9364 14746 9430 14756
rect 9556 14746 9622 14756
rect 9748 14746 9814 14756
rect 9940 14746 10006 14756
rect 10132 14746 10198 14756
rect 10324 14746 10390 14756
rect 10516 14746 10582 14756
rect 11000 14746 11066 14756
rect 11192 14746 11258 14756
rect 11384 14746 11450 14756
rect 11576 14746 11642 14756
rect 11768 14746 11834 14756
rect 11960 14746 12026 14756
rect 12152 14746 12218 14756
rect 12344 14746 12410 14756
rect 12828 14746 12894 14756
rect 13020 14746 13086 14756
rect 13212 14746 13278 14756
rect 13404 14746 13470 14756
rect 13596 14746 13662 14756
rect 13788 14746 13854 14756
rect 13980 14746 14046 14756
rect 14172 14746 14238 14756
rect 14656 14746 14722 14756
rect 14848 14746 14914 14756
rect 15040 14746 15106 14756
rect 15232 14746 15298 14756
rect 15424 14746 15490 14756
rect 15616 14746 15682 14756
rect 15808 14746 15874 14756
rect 16000 14746 16066 14756
rect 16484 14746 16550 14756
rect 16676 14746 16742 14756
rect 16868 14746 16934 14756
rect 17060 14746 17126 14756
rect 17252 14746 17318 14756
rect 17444 14746 17510 14756
rect 17636 14746 17702 14756
rect 17828 14746 17894 14756
rect 18312 14746 18378 14756
rect 18504 14746 18570 14756
rect 18696 14746 18762 14756
rect 18888 14746 18954 14756
rect 19080 14746 19146 14756
rect 19272 14746 19338 14756
rect 19464 14746 19530 14756
rect 19656 14746 19722 14756
rect 20140 14746 20206 14756
rect 20332 14746 20398 14756
rect 20524 14746 20590 14756
rect 20716 14746 20782 14756
rect 20908 14746 20974 14756
rect 21100 14746 21166 14756
rect 21292 14746 21358 14756
rect 21484 14746 21550 14756
rect 0 14593 32 14746
rect 98 14593 224 14746
rect 290 14593 416 14746
rect 482 14593 608 14746
rect 674 14593 800 14746
rect 866 14593 992 14746
rect 1058 14593 1184 14746
rect 1250 14593 1376 14746
rect 1828 14593 1860 14746
rect 1926 14593 2052 14746
rect 2118 14593 2244 14746
rect 2310 14593 2436 14746
rect 2502 14593 2628 14746
rect 2694 14593 2820 14746
rect 2886 14593 3012 14746
rect 3078 14593 3204 14746
rect 3656 14593 3688 14746
rect 3754 14593 3880 14746
rect 3946 14593 4072 14746
rect 4138 14593 4264 14746
rect 4330 14593 4456 14746
rect 4522 14593 4648 14746
rect 4714 14593 4840 14746
rect 4906 14593 5032 14746
rect 5484 14593 5516 14746
rect 5582 14593 5708 14746
rect 5774 14593 5900 14746
rect 5966 14593 6092 14746
rect 6158 14593 6284 14746
rect 6350 14593 6476 14746
rect 6542 14593 6668 14746
rect 6734 14593 6860 14746
rect 7312 14593 7344 14746
rect 7410 14593 7536 14746
rect 7602 14593 7728 14746
rect 7794 14593 7920 14746
rect 7986 14593 8112 14746
rect 8178 14593 8304 14746
rect 8370 14593 8496 14746
rect 8562 14593 8688 14746
rect 9140 14593 9172 14746
rect 9238 14593 9364 14746
rect 9430 14593 9556 14746
rect 9622 14593 9748 14746
rect 9814 14593 9940 14746
rect 10006 14593 10132 14746
rect 10198 14593 10324 14746
rect 10390 14593 10516 14746
rect 10968 14593 11000 14746
rect 11066 14593 11192 14746
rect 11258 14593 11384 14746
rect 11450 14593 11576 14746
rect 11642 14593 11768 14746
rect 11834 14593 11960 14746
rect 12026 14593 12152 14746
rect 12218 14593 12344 14746
rect 12796 14593 12828 14746
rect 12894 14593 13020 14746
rect 13086 14593 13212 14746
rect 13278 14593 13404 14746
rect 13470 14593 13596 14746
rect 13662 14593 13788 14746
rect 13854 14593 13980 14746
rect 14046 14593 14172 14746
rect 14624 14593 14656 14746
rect 14722 14593 14848 14746
rect 14914 14593 15040 14746
rect 15106 14593 15232 14746
rect 15298 14593 15424 14746
rect 15490 14593 15616 14746
rect 15682 14593 15808 14746
rect 15874 14593 16000 14746
rect 16452 14593 16484 14746
rect 16550 14593 16676 14746
rect 16742 14593 16868 14746
rect 16934 14593 17060 14746
rect 17126 14593 17252 14746
rect 17318 14593 17444 14746
rect 17510 14593 17636 14746
rect 17702 14593 17828 14746
rect 18280 14593 18312 14746
rect 18378 14593 18504 14746
rect 18570 14593 18696 14746
rect 18762 14593 18888 14746
rect 18954 14593 19080 14746
rect 19146 14593 19272 14746
rect 19338 14593 19464 14746
rect 19530 14593 19656 14746
rect 20108 14593 20140 14746
rect 20206 14593 20332 14746
rect 20398 14593 20524 14746
rect 20590 14593 20716 14746
rect 20782 14593 20908 14746
rect 20974 14593 21100 14746
rect 21166 14593 21292 14746
rect 21358 14593 21484 14746
rect 32 14583 98 14593
rect 224 14583 290 14593
rect 416 14583 482 14593
rect 608 14583 674 14593
rect 800 14583 866 14593
rect 992 14583 1058 14593
rect 1184 14583 1250 14593
rect 1376 14583 1442 14593
rect 1860 14583 1926 14593
rect 2052 14583 2118 14593
rect 2244 14583 2310 14593
rect 2436 14583 2502 14593
rect 2628 14583 2694 14593
rect 2820 14583 2886 14593
rect 3012 14583 3078 14593
rect 3204 14583 3270 14593
rect 3688 14583 3754 14593
rect 3880 14583 3946 14593
rect 4072 14583 4138 14593
rect 4264 14583 4330 14593
rect 4456 14583 4522 14593
rect 4648 14583 4714 14593
rect 4840 14583 4906 14593
rect 5032 14583 5098 14593
rect 5516 14583 5582 14593
rect 5708 14583 5774 14593
rect 5900 14583 5966 14593
rect 6092 14583 6158 14593
rect 6284 14583 6350 14593
rect 6476 14583 6542 14593
rect 6668 14583 6734 14593
rect 6860 14583 6926 14593
rect 7344 14583 7410 14593
rect 7536 14583 7602 14593
rect 7728 14583 7794 14593
rect 7920 14583 7986 14593
rect 8112 14583 8178 14593
rect 8304 14583 8370 14593
rect 8496 14583 8562 14593
rect 8688 14583 8754 14593
rect 9172 14583 9238 14593
rect 9364 14583 9430 14593
rect 9556 14583 9622 14593
rect 9748 14583 9814 14593
rect 9940 14583 10006 14593
rect 10132 14583 10198 14593
rect 10324 14583 10390 14593
rect 10516 14583 10582 14593
rect 11000 14583 11066 14593
rect 11192 14583 11258 14593
rect 11384 14583 11450 14593
rect 11576 14583 11642 14593
rect 11768 14583 11834 14593
rect 11960 14583 12026 14593
rect 12152 14583 12218 14593
rect 12344 14583 12410 14593
rect 12828 14583 12894 14593
rect 13020 14583 13086 14593
rect 13212 14583 13278 14593
rect 13404 14583 13470 14593
rect 13596 14583 13662 14593
rect 13788 14583 13854 14593
rect 13980 14583 14046 14593
rect 14172 14583 14238 14593
rect 14656 14583 14722 14593
rect 14848 14583 14914 14593
rect 15040 14583 15106 14593
rect 15232 14583 15298 14593
rect 15424 14583 15490 14593
rect 15616 14583 15682 14593
rect 15808 14583 15874 14593
rect 16000 14583 16066 14593
rect 16484 14583 16550 14593
rect 16676 14583 16742 14593
rect 16868 14583 16934 14593
rect 17060 14583 17126 14593
rect 17252 14583 17318 14593
rect 17444 14583 17510 14593
rect 17636 14583 17702 14593
rect 17828 14583 17894 14593
rect 18312 14583 18378 14593
rect 18504 14583 18570 14593
rect 18696 14583 18762 14593
rect 18888 14583 18954 14593
rect 19080 14583 19146 14593
rect 19272 14583 19338 14593
rect 19464 14583 19530 14593
rect 19656 14583 19722 14593
rect 20140 14583 20206 14593
rect 20332 14583 20398 14593
rect 20524 14583 20590 14593
rect 20716 14583 20782 14593
rect 20908 14583 20974 14593
rect 21100 14583 21166 14593
rect 21292 14583 21358 14593
rect 21484 14583 21550 14593
rect 128 14533 194 14543
rect 320 14533 386 14543
rect 512 14533 578 14543
rect 704 14533 770 14543
rect 896 14533 962 14543
rect 1088 14533 1154 14543
rect 1280 14533 1346 14543
rect 1472 14533 1528 14543
rect 1956 14533 2022 14543
rect 2148 14533 2214 14543
rect 2340 14533 2406 14543
rect 2532 14533 2598 14543
rect 2724 14533 2790 14543
rect 2916 14533 2982 14543
rect 3108 14533 3174 14543
rect 3300 14533 3356 14543
rect 3784 14533 3850 14543
rect 3976 14533 4042 14543
rect 4168 14533 4234 14543
rect 4360 14533 4426 14543
rect 4552 14533 4618 14543
rect 4744 14533 4810 14543
rect 4936 14533 5002 14543
rect 5128 14533 5184 14543
rect 5612 14533 5678 14543
rect 5804 14533 5870 14543
rect 5996 14533 6062 14543
rect 6188 14533 6254 14543
rect 6380 14533 6446 14543
rect 6572 14533 6638 14543
rect 6764 14533 6830 14543
rect 6956 14533 7012 14543
rect 7440 14533 7506 14543
rect 7632 14533 7698 14543
rect 7824 14533 7890 14543
rect 8016 14533 8082 14543
rect 8208 14533 8274 14543
rect 8400 14533 8466 14543
rect 8592 14533 8658 14543
rect 8784 14533 8840 14543
rect 9268 14533 9334 14543
rect 9460 14533 9526 14543
rect 9652 14533 9718 14543
rect 9844 14533 9910 14543
rect 10036 14533 10102 14543
rect 10228 14533 10294 14543
rect 10420 14533 10486 14543
rect 10612 14533 10668 14543
rect 11096 14533 11162 14543
rect 11288 14533 11354 14543
rect 11480 14533 11546 14543
rect 11672 14533 11738 14543
rect 11864 14533 11930 14543
rect 12056 14533 12122 14543
rect 12248 14533 12314 14543
rect 12440 14533 12496 14543
rect 12924 14533 12990 14543
rect 13116 14533 13182 14543
rect 13308 14533 13374 14543
rect 13500 14533 13566 14543
rect 13692 14533 13758 14543
rect 13884 14533 13950 14543
rect 14076 14533 14142 14543
rect 14268 14533 14324 14543
rect 14752 14533 14818 14543
rect 14944 14533 15010 14543
rect 15136 14533 15202 14543
rect 15328 14533 15394 14543
rect 15520 14533 15586 14543
rect 15712 14533 15778 14543
rect 15904 14533 15970 14543
rect 16096 14533 16152 14543
rect 16580 14533 16646 14543
rect 16772 14533 16838 14543
rect 16964 14533 17030 14543
rect 17156 14533 17222 14543
rect 17348 14533 17414 14543
rect 17540 14533 17606 14543
rect 17732 14533 17798 14543
rect 17924 14533 17980 14543
rect 18408 14533 18474 14543
rect 18600 14533 18666 14543
rect 18792 14533 18858 14543
rect 18984 14533 19050 14543
rect 19176 14533 19242 14543
rect 19368 14533 19434 14543
rect 19560 14533 19626 14543
rect 19752 14533 19808 14543
rect 20236 14533 20302 14543
rect 20428 14533 20494 14543
rect 20620 14533 20686 14543
rect 20812 14533 20878 14543
rect 21004 14533 21070 14543
rect 21196 14533 21262 14543
rect 21388 14533 21454 14543
rect 21580 14533 21636 14543
rect 0 14380 128 14533
rect 194 14380 320 14533
rect 386 14380 512 14533
rect 578 14380 704 14533
rect 770 14380 896 14533
rect 962 14380 1088 14533
rect 1154 14380 1280 14533
rect 1346 14380 1472 14533
rect 1528 14380 1708 14533
rect 1828 14380 1956 14533
rect 2022 14380 2148 14533
rect 2214 14380 2340 14533
rect 2406 14380 2532 14533
rect 2598 14380 2724 14533
rect 2790 14380 2916 14533
rect 2982 14380 3108 14533
rect 3174 14380 3300 14533
rect 3356 14380 3536 14533
rect 3656 14380 3784 14533
rect 3850 14380 3976 14533
rect 4042 14380 4168 14533
rect 4234 14380 4360 14533
rect 4426 14380 4552 14533
rect 4618 14380 4744 14533
rect 4810 14380 4936 14533
rect 5002 14380 5128 14533
rect 5184 14380 5364 14533
rect 5484 14380 5612 14533
rect 5678 14380 5804 14533
rect 5870 14380 5996 14533
rect 6062 14380 6188 14533
rect 6254 14380 6380 14533
rect 6446 14380 6572 14533
rect 6638 14380 6764 14533
rect 6830 14380 6956 14533
rect 7012 14380 7192 14533
rect 7312 14380 7440 14533
rect 7506 14380 7632 14533
rect 7698 14380 7824 14533
rect 7890 14380 8016 14533
rect 8082 14380 8208 14533
rect 8274 14380 8400 14533
rect 8466 14380 8592 14533
rect 8658 14380 8784 14533
rect 8840 14380 9020 14533
rect 9140 14380 9268 14533
rect 9334 14380 9460 14533
rect 9526 14380 9652 14533
rect 9718 14380 9844 14533
rect 9910 14380 10036 14533
rect 10102 14380 10228 14533
rect 10294 14380 10420 14533
rect 10486 14380 10612 14533
rect 10668 14380 10848 14533
rect 10968 14380 11096 14533
rect 11162 14380 11288 14533
rect 11354 14380 11480 14533
rect 11546 14380 11672 14533
rect 11738 14380 11864 14533
rect 11930 14380 12056 14533
rect 12122 14380 12248 14533
rect 12314 14380 12440 14533
rect 12496 14380 12676 14533
rect 12796 14380 12924 14533
rect 12990 14380 13116 14533
rect 13182 14380 13308 14533
rect 13374 14380 13500 14533
rect 13566 14380 13692 14533
rect 13758 14380 13884 14533
rect 13950 14380 14076 14533
rect 14142 14380 14268 14533
rect 14324 14380 14504 14533
rect 14624 14380 14752 14533
rect 14818 14380 14944 14533
rect 15010 14380 15136 14533
rect 15202 14380 15328 14533
rect 15394 14380 15520 14533
rect 15586 14380 15712 14533
rect 15778 14380 15904 14533
rect 15970 14380 16096 14533
rect 16152 14380 16332 14533
rect 16452 14380 16580 14533
rect 16646 14380 16772 14533
rect 16838 14380 16964 14533
rect 17030 14380 17156 14533
rect 17222 14380 17348 14533
rect 17414 14380 17540 14533
rect 17606 14380 17732 14533
rect 17798 14380 17924 14533
rect 17980 14380 18160 14533
rect 18280 14380 18408 14533
rect 18474 14380 18600 14533
rect 18666 14380 18792 14533
rect 18858 14380 18984 14533
rect 19050 14380 19176 14533
rect 19242 14380 19368 14533
rect 19434 14380 19560 14533
rect 19626 14380 19752 14533
rect 19808 14380 19988 14533
rect 20108 14380 20236 14533
rect 20302 14380 20428 14533
rect 20494 14380 20620 14533
rect 20686 14380 20812 14533
rect 20878 14380 21004 14533
rect 21070 14380 21196 14533
rect 21262 14380 21388 14533
rect 21454 14380 21580 14533
rect 21636 14380 21816 14533
rect 128 14370 194 14380
rect 320 14370 386 14380
rect 512 14370 578 14380
rect 704 14370 770 14380
rect 896 14370 962 14380
rect 1088 14370 1154 14380
rect 1280 14370 1346 14380
rect 1472 14370 1528 14380
rect 1956 14370 2022 14380
rect 2148 14370 2214 14380
rect 2340 14370 2406 14380
rect 2532 14370 2598 14380
rect 2724 14370 2790 14380
rect 2916 14370 2982 14380
rect 3108 14370 3174 14380
rect 3300 14370 3356 14380
rect 3784 14370 3850 14380
rect 3976 14370 4042 14380
rect 4168 14370 4234 14380
rect 4360 14370 4426 14380
rect 4552 14370 4618 14380
rect 4744 14370 4810 14380
rect 4936 14370 5002 14380
rect 5128 14370 5184 14380
rect 5612 14370 5678 14380
rect 5804 14370 5870 14380
rect 5996 14370 6062 14380
rect 6188 14370 6254 14380
rect 6380 14370 6446 14380
rect 6572 14370 6638 14380
rect 6764 14370 6830 14380
rect 6956 14370 7012 14380
rect 7440 14370 7506 14380
rect 7632 14370 7698 14380
rect 7824 14370 7890 14380
rect 8016 14370 8082 14380
rect 8208 14370 8274 14380
rect 8400 14370 8466 14380
rect 8592 14370 8658 14380
rect 8784 14370 8840 14380
rect 9268 14370 9334 14380
rect 9460 14370 9526 14380
rect 9652 14370 9718 14380
rect 9844 14370 9910 14380
rect 10036 14370 10102 14380
rect 10228 14370 10294 14380
rect 10420 14370 10486 14380
rect 10612 14370 10668 14380
rect 11096 14370 11162 14380
rect 11288 14370 11354 14380
rect 11480 14370 11546 14380
rect 11672 14370 11738 14380
rect 11864 14370 11930 14380
rect 12056 14370 12122 14380
rect 12248 14370 12314 14380
rect 12440 14370 12496 14380
rect 12924 14370 12990 14380
rect 13116 14370 13182 14380
rect 13308 14370 13374 14380
rect 13500 14370 13566 14380
rect 13692 14370 13758 14380
rect 13884 14370 13950 14380
rect 14076 14370 14142 14380
rect 14268 14370 14324 14380
rect 14752 14370 14818 14380
rect 14944 14370 15010 14380
rect 15136 14370 15202 14380
rect 15328 14370 15394 14380
rect 15520 14370 15586 14380
rect 15712 14370 15778 14380
rect 15904 14370 15970 14380
rect 16096 14370 16152 14380
rect 16580 14370 16646 14380
rect 16772 14370 16838 14380
rect 16964 14370 17030 14380
rect 17156 14370 17222 14380
rect 17348 14370 17414 14380
rect 17540 14370 17606 14380
rect 17732 14370 17798 14380
rect 17924 14370 17980 14380
rect 18408 14370 18474 14380
rect 18600 14370 18666 14380
rect 18792 14370 18858 14380
rect 18984 14370 19050 14380
rect 19176 14370 19242 14380
rect 19368 14370 19434 14380
rect 19560 14370 19626 14380
rect 19752 14370 19808 14380
rect 20236 14370 20302 14380
rect 20428 14370 20494 14380
rect 20620 14370 20686 14380
rect 20812 14370 20878 14380
rect 21004 14370 21070 14380
rect 21196 14370 21262 14380
rect 21388 14370 21454 14380
rect 21580 14370 21636 14380
rect 32 14032 98 14042
rect 224 14032 290 14042
rect 416 14032 482 14042
rect 608 14032 674 14042
rect 800 14032 866 14042
rect 992 14032 1058 14042
rect 1184 14032 1250 14042
rect 1376 14032 1442 14042
rect 1860 14032 1926 14042
rect 2052 14032 2118 14042
rect 2244 14032 2310 14042
rect 2436 14032 2502 14042
rect 2628 14032 2694 14042
rect 2820 14032 2886 14042
rect 3012 14032 3078 14042
rect 3204 14032 3270 14042
rect 3688 14032 3754 14042
rect 3880 14032 3946 14042
rect 4072 14032 4138 14042
rect 4264 14032 4330 14042
rect 4456 14032 4522 14042
rect 4648 14032 4714 14042
rect 4840 14032 4906 14042
rect 5032 14032 5098 14042
rect 5516 14032 5582 14042
rect 5708 14032 5774 14042
rect 5900 14032 5966 14042
rect 6092 14032 6158 14042
rect 6284 14032 6350 14042
rect 6476 14032 6542 14042
rect 6668 14032 6734 14042
rect 6860 14032 6926 14042
rect 7344 14032 7410 14042
rect 7536 14032 7602 14042
rect 7728 14032 7794 14042
rect 7920 14032 7986 14042
rect 8112 14032 8178 14042
rect 8304 14032 8370 14042
rect 8496 14032 8562 14042
rect 8688 14032 8754 14042
rect 9172 14032 9238 14042
rect 9364 14032 9430 14042
rect 9556 14032 9622 14042
rect 9748 14032 9814 14042
rect 9940 14032 10006 14042
rect 10132 14032 10198 14042
rect 10324 14032 10390 14042
rect 10516 14032 10582 14042
rect 11000 14032 11066 14042
rect 11192 14032 11258 14042
rect 11384 14032 11450 14042
rect 11576 14032 11642 14042
rect 11768 14032 11834 14042
rect 11960 14032 12026 14042
rect 12152 14032 12218 14042
rect 12344 14032 12410 14042
rect 12828 14032 12894 14042
rect 13020 14032 13086 14042
rect 13212 14032 13278 14042
rect 13404 14032 13470 14042
rect 13596 14032 13662 14042
rect 13788 14032 13854 14042
rect 13980 14032 14046 14042
rect 14172 14032 14238 14042
rect 14656 14032 14722 14042
rect 14848 14032 14914 14042
rect 15040 14032 15106 14042
rect 15232 14032 15298 14042
rect 15424 14032 15490 14042
rect 15616 14032 15682 14042
rect 15808 14032 15874 14042
rect 16000 14032 16066 14042
rect 16484 14032 16550 14042
rect 16676 14032 16742 14042
rect 16868 14032 16934 14042
rect 17060 14032 17126 14042
rect 17252 14032 17318 14042
rect 17444 14032 17510 14042
rect 17636 14032 17702 14042
rect 17828 14032 17894 14042
rect 18312 14032 18378 14042
rect 18504 14032 18570 14042
rect 18696 14032 18762 14042
rect 18888 14032 18954 14042
rect 19080 14032 19146 14042
rect 19272 14032 19338 14042
rect 19464 14032 19530 14042
rect 19656 14032 19722 14042
rect 20140 14032 20206 14042
rect 20332 14032 20398 14042
rect 20524 14032 20590 14042
rect 20716 14032 20782 14042
rect 20908 14032 20974 14042
rect 21100 14032 21166 14042
rect 21292 14032 21358 14042
rect 21484 14032 21550 14042
rect 0 13879 32 14032
rect 98 13879 224 14032
rect 290 13879 416 14032
rect 482 13879 608 14032
rect 674 13879 800 14032
rect 866 13879 992 14032
rect 1058 13879 1184 14032
rect 1250 13879 1376 14032
rect 1828 13879 1860 14032
rect 1926 13879 2052 14032
rect 2118 13879 2244 14032
rect 2310 13879 2436 14032
rect 2502 13879 2628 14032
rect 2694 13879 2820 14032
rect 2886 13879 3012 14032
rect 3078 13879 3204 14032
rect 3656 13879 3688 14032
rect 3754 13879 3880 14032
rect 3946 13879 4072 14032
rect 4138 13879 4264 14032
rect 4330 13879 4456 14032
rect 4522 13879 4648 14032
rect 4714 13879 4840 14032
rect 4906 13879 5032 14032
rect 5484 13879 5516 14032
rect 5582 13879 5708 14032
rect 5774 13879 5900 14032
rect 5966 13879 6092 14032
rect 6158 13879 6284 14032
rect 6350 13879 6476 14032
rect 6542 13879 6668 14032
rect 6734 13879 6860 14032
rect 7312 13879 7344 14032
rect 7410 13879 7536 14032
rect 7602 13879 7728 14032
rect 7794 13879 7920 14032
rect 7986 13879 8112 14032
rect 8178 13879 8304 14032
rect 8370 13879 8496 14032
rect 8562 13879 8688 14032
rect 9140 13879 9172 14032
rect 9238 13879 9364 14032
rect 9430 13879 9556 14032
rect 9622 13879 9748 14032
rect 9814 13879 9940 14032
rect 10006 13879 10132 14032
rect 10198 13879 10324 14032
rect 10390 13879 10516 14032
rect 10968 13879 11000 14032
rect 11066 13879 11192 14032
rect 11258 13879 11384 14032
rect 11450 13879 11576 14032
rect 11642 13879 11768 14032
rect 11834 13879 11960 14032
rect 12026 13879 12152 14032
rect 12218 13879 12344 14032
rect 12796 13879 12828 14032
rect 12894 13879 13020 14032
rect 13086 13879 13212 14032
rect 13278 13879 13404 14032
rect 13470 13879 13596 14032
rect 13662 13879 13788 14032
rect 13854 13879 13980 14032
rect 14046 13879 14172 14032
rect 14624 13879 14656 14032
rect 14722 13879 14848 14032
rect 14914 13879 15040 14032
rect 15106 13879 15232 14032
rect 15298 13879 15424 14032
rect 15490 13879 15616 14032
rect 15682 13879 15808 14032
rect 15874 13879 16000 14032
rect 16452 13879 16484 14032
rect 16550 13879 16676 14032
rect 16742 13879 16868 14032
rect 16934 13879 17060 14032
rect 17126 13879 17252 14032
rect 17318 13879 17444 14032
rect 17510 13879 17636 14032
rect 17702 13879 17828 14032
rect 18280 13879 18312 14032
rect 18378 13879 18504 14032
rect 18570 13879 18696 14032
rect 18762 13879 18888 14032
rect 18954 13879 19080 14032
rect 19146 13879 19272 14032
rect 19338 13879 19464 14032
rect 19530 13879 19656 14032
rect 20108 13879 20140 14032
rect 20206 13879 20332 14032
rect 20398 13879 20524 14032
rect 20590 13879 20716 14032
rect 20782 13879 20908 14032
rect 20974 13879 21100 14032
rect 21166 13879 21292 14032
rect 21358 13879 21484 14032
rect 32 13869 98 13879
rect 224 13869 290 13879
rect 416 13869 482 13879
rect 608 13869 674 13879
rect 800 13869 866 13879
rect 992 13869 1058 13879
rect 1184 13869 1250 13879
rect 1376 13869 1442 13879
rect 1860 13869 1926 13879
rect 2052 13869 2118 13879
rect 2244 13869 2310 13879
rect 2436 13869 2502 13879
rect 2628 13869 2694 13879
rect 2820 13869 2886 13879
rect 3012 13869 3078 13879
rect 3204 13869 3270 13879
rect 3688 13869 3754 13879
rect 3880 13869 3946 13879
rect 4072 13869 4138 13879
rect 4264 13869 4330 13879
rect 4456 13869 4522 13879
rect 4648 13869 4714 13879
rect 4840 13869 4906 13879
rect 5032 13869 5098 13879
rect 5516 13869 5582 13879
rect 5708 13869 5774 13879
rect 5900 13869 5966 13879
rect 6092 13869 6158 13879
rect 6284 13869 6350 13879
rect 6476 13869 6542 13879
rect 6668 13869 6734 13879
rect 6860 13869 6926 13879
rect 7344 13869 7410 13879
rect 7536 13869 7602 13879
rect 7728 13869 7794 13879
rect 7920 13869 7986 13879
rect 8112 13869 8178 13879
rect 8304 13869 8370 13879
rect 8496 13869 8562 13879
rect 8688 13869 8754 13879
rect 9172 13869 9238 13879
rect 9364 13869 9430 13879
rect 9556 13869 9622 13879
rect 9748 13869 9814 13879
rect 9940 13869 10006 13879
rect 10132 13869 10198 13879
rect 10324 13869 10390 13879
rect 10516 13869 10582 13879
rect 11000 13869 11066 13879
rect 11192 13869 11258 13879
rect 11384 13869 11450 13879
rect 11576 13869 11642 13879
rect 11768 13869 11834 13879
rect 11960 13869 12026 13879
rect 12152 13869 12218 13879
rect 12344 13869 12410 13879
rect 12828 13869 12894 13879
rect 13020 13869 13086 13879
rect 13212 13869 13278 13879
rect 13404 13869 13470 13879
rect 13596 13869 13662 13879
rect 13788 13869 13854 13879
rect 13980 13869 14046 13879
rect 14172 13869 14238 13879
rect 14656 13869 14722 13879
rect 14848 13869 14914 13879
rect 15040 13869 15106 13879
rect 15232 13869 15298 13879
rect 15424 13869 15490 13879
rect 15616 13869 15682 13879
rect 15808 13869 15874 13879
rect 16000 13869 16066 13879
rect 16484 13869 16550 13879
rect 16676 13869 16742 13879
rect 16868 13869 16934 13879
rect 17060 13869 17126 13879
rect 17252 13869 17318 13879
rect 17444 13869 17510 13879
rect 17636 13869 17702 13879
rect 17828 13869 17894 13879
rect 18312 13869 18378 13879
rect 18504 13869 18570 13879
rect 18696 13869 18762 13879
rect 18888 13869 18954 13879
rect 19080 13869 19146 13879
rect 19272 13869 19338 13879
rect 19464 13869 19530 13879
rect 19656 13869 19722 13879
rect 20140 13869 20206 13879
rect 20332 13869 20398 13879
rect 20524 13869 20590 13879
rect 20716 13869 20782 13879
rect 20908 13869 20974 13879
rect 21100 13869 21166 13879
rect 21292 13869 21358 13879
rect 21484 13869 21550 13879
rect 128 13819 194 13829
rect 320 13819 386 13829
rect 512 13819 578 13829
rect 704 13819 770 13829
rect 896 13819 962 13829
rect 1088 13819 1154 13829
rect 1280 13819 1346 13829
rect 1472 13819 1528 13829
rect 1956 13819 2022 13829
rect 2148 13819 2214 13829
rect 2340 13819 2406 13829
rect 2532 13819 2598 13829
rect 2724 13819 2790 13829
rect 2916 13819 2982 13829
rect 3108 13819 3174 13829
rect 3300 13819 3356 13829
rect 3784 13819 3850 13829
rect 3976 13819 4042 13829
rect 4168 13819 4234 13829
rect 4360 13819 4426 13829
rect 4552 13819 4618 13829
rect 4744 13819 4810 13829
rect 4936 13819 5002 13829
rect 5128 13819 5184 13829
rect 5612 13819 5678 13829
rect 5804 13819 5870 13829
rect 5996 13819 6062 13829
rect 6188 13819 6254 13829
rect 6380 13819 6446 13829
rect 6572 13819 6638 13829
rect 6764 13819 6830 13829
rect 6956 13819 7012 13829
rect 7440 13819 7506 13829
rect 7632 13819 7698 13829
rect 7824 13819 7890 13829
rect 8016 13819 8082 13829
rect 8208 13819 8274 13829
rect 8400 13819 8466 13829
rect 8592 13819 8658 13829
rect 8784 13819 8840 13829
rect 9268 13819 9334 13829
rect 9460 13819 9526 13829
rect 9652 13819 9718 13829
rect 9844 13819 9910 13829
rect 10036 13819 10102 13829
rect 10228 13819 10294 13829
rect 10420 13819 10486 13829
rect 10612 13819 10668 13829
rect 11096 13819 11162 13829
rect 11288 13819 11354 13829
rect 11480 13819 11546 13829
rect 11672 13819 11738 13829
rect 11864 13819 11930 13829
rect 12056 13819 12122 13829
rect 12248 13819 12314 13829
rect 12440 13819 12496 13829
rect 12924 13819 12990 13829
rect 13116 13819 13182 13829
rect 13308 13819 13374 13829
rect 13500 13819 13566 13829
rect 13692 13819 13758 13829
rect 13884 13819 13950 13829
rect 14076 13819 14142 13829
rect 14268 13819 14324 13829
rect 14752 13819 14818 13829
rect 14944 13819 15010 13829
rect 15136 13819 15202 13829
rect 15328 13819 15394 13829
rect 15520 13819 15586 13829
rect 15712 13819 15778 13829
rect 15904 13819 15970 13829
rect 16096 13819 16152 13829
rect 16580 13819 16646 13829
rect 16772 13819 16838 13829
rect 16964 13819 17030 13829
rect 17156 13819 17222 13829
rect 17348 13819 17414 13829
rect 17540 13819 17606 13829
rect 17732 13819 17798 13829
rect 17924 13819 17980 13829
rect 18408 13819 18474 13829
rect 18600 13819 18666 13829
rect 18792 13819 18858 13829
rect 18984 13819 19050 13829
rect 19176 13819 19242 13829
rect 19368 13819 19434 13829
rect 19560 13819 19626 13829
rect 19752 13819 19808 13829
rect 20236 13819 20302 13829
rect 20428 13819 20494 13829
rect 20620 13819 20686 13829
rect 20812 13819 20878 13829
rect 21004 13819 21070 13829
rect 21196 13819 21262 13829
rect 21388 13819 21454 13829
rect 21580 13819 21636 13829
rect 0 13666 128 13819
rect 194 13666 320 13819
rect 386 13666 512 13819
rect 578 13666 704 13819
rect 770 13666 896 13819
rect 962 13666 1088 13819
rect 1154 13666 1280 13819
rect 1346 13666 1472 13819
rect 1528 13666 1708 13819
rect 1828 13666 1956 13819
rect 2022 13666 2148 13819
rect 2214 13666 2340 13819
rect 2406 13666 2532 13819
rect 2598 13666 2724 13819
rect 2790 13666 2916 13819
rect 2982 13666 3108 13819
rect 3174 13666 3300 13819
rect 3356 13666 3536 13819
rect 3656 13666 3784 13819
rect 3850 13666 3976 13819
rect 4042 13666 4168 13819
rect 4234 13666 4360 13819
rect 4426 13666 4552 13819
rect 4618 13666 4744 13819
rect 4810 13666 4936 13819
rect 5002 13666 5128 13819
rect 5184 13666 5364 13819
rect 5484 13666 5612 13819
rect 5678 13666 5804 13819
rect 5870 13666 5996 13819
rect 6062 13666 6188 13819
rect 6254 13666 6380 13819
rect 6446 13666 6572 13819
rect 6638 13666 6764 13819
rect 6830 13666 6956 13819
rect 7012 13666 7192 13819
rect 7312 13666 7440 13819
rect 7506 13666 7632 13819
rect 7698 13666 7824 13819
rect 7890 13666 8016 13819
rect 8082 13666 8208 13819
rect 8274 13666 8400 13819
rect 8466 13666 8592 13819
rect 8658 13666 8784 13819
rect 8840 13666 9020 13819
rect 9140 13666 9268 13819
rect 9334 13666 9460 13819
rect 9526 13666 9652 13819
rect 9718 13666 9844 13819
rect 9910 13666 10036 13819
rect 10102 13666 10228 13819
rect 10294 13666 10420 13819
rect 10486 13666 10612 13819
rect 10668 13666 10848 13819
rect 10968 13666 11096 13819
rect 11162 13666 11288 13819
rect 11354 13666 11480 13819
rect 11546 13666 11672 13819
rect 11738 13666 11864 13819
rect 11930 13666 12056 13819
rect 12122 13666 12248 13819
rect 12314 13666 12440 13819
rect 12496 13666 12676 13819
rect 12796 13666 12924 13819
rect 12990 13666 13116 13819
rect 13182 13666 13308 13819
rect 13374 13666 13500 13819
rect 13566 13666 13692 13819
rect 13758 13666 13884 13819
rect 13950 13666 14076 13819
rect 14142 13666 14268 13819
rect 14324 13666 14504 13819
rect 14624 13666 14752 13819
rect 14818 13666 14944 13819
rect 15010 13666 15136 13819
rect 15202 13666 15328 13819
rect 15394 13666 15520 13819
rect 15586 13666 15712 13819
rect 15778 13666 15904 13819
rect 15970 13666 16096 13819
rect 16152 13666 16332 13819
rect 16452 13666 16580 13819
rect 16646 13666 16772 13819
rect 16838 13666 16964 13819
rect 17030 13666 17156 13819
rect 17222 13666 17348 13819
rect 17414 13666 17540 13819
rect 17606 13666 17732 13819
rect 17798 13666 17924 13819
rect 17980 13666 18160 13819
rect 18280 13666 18408 13819
rect 18474 13666 18600 13819
rect 18666 13666 18792 13819
rect 18858 13666 18984 13819
rect 19050 13666 19176 13819
rect 19242 13666 19368 13819
rect 19434 13666 19560 13819
rect 19626 13666 19752 13819
rect 19808 13666 19988 13819
rect 20108 13666 20236 13819
rect 20302 13666 20428 13819
rect 20494 13666 20620 13819
rect 20686 13666 20812 13819
rect 20878 13666 21004 13819
rect 21070 13666 21196 13819
rect 21262 13666 21388 13819
rect 21454 13666 21580 13819
rect 21636 13666 21816 13819
rect 128 13656 194 13666
rect 320 13656 386 13666
rect 512 13656 578 13666
rect 704 13656 770 13666
rect 896 13656 962 13666
rect 1088 13656 1154 13666
rect 1280 13656 1346 13666
rect 1472 13656 1528 13666
rect 1956 13656 2022 13666
rect 2148 13656 2214 13666
rect 2340 13656 2406 13666
rect 2532 13656 2598 13666
rect 2724 13656 2790 13666
rect 2916 13656 2982 13666
rect 3108 13656 3174 13666
rect 3300 13656 3356 13666
rect 3784 13656 3850 13666
rect 3976 13656 4042 13666
rect 4168 13656 4234 13666
rect 4360 13656 4426 13666
rect 4552 13656 4618 13666
rect 4744 13656 4810 13666
rect 4936 13656 5002 13666
rect 5128 13656 5184 13666
rect 5612 13656 5678 13666
rect 5804 13656 5870 13666
rect 5996 13656 6062 13666
rect 6188 13656 6254 13666
rect 6380 13656 6446 13666
rect 6572 13656 6638 13666
rect 6764 13656 6830 13666
rect 6956 13656 7012 13666
rect 7440 13656 7506 13666
rect 7632 13656 7698 13666
rect 7824 13656 7890 13666
rect 8016 13656 8082 13666
rect 8208 13656 8274 13666
rect 8400 13656 8466 13666
rect 8592 13656 8658 13666
rect 8784 13656 8840 13666
rect 9268 13656 9334 13666
rect 9460 13656 9526 13666
rect 9652 13656 9718 13666
rect 9844 13656 9910 13666
rect 10036 13656 10102 13666
rect 10228 13656 10294 13666
rect 10420 13656 10486 13666
rect 10612 13656 10668 13666
rect 11096 13656 11162 13666
rect 11288 13656 11354 13666
rect 11480 13656 11546 13666
rect 11672 13656 11738 13666
rect 11864 13656 11930 13666
rect 12056 13656 12122 13666
rect 12248 13656 12314 13666
rect 12440 13656 12496 13666
rect 12924 13656 12990 13666
rect 13116 13656 13182 13666
rect 13308 13656 13374 13666
rect 13500 13656 13566 13666
rect 13692 13656 13758 13666
rect 13884 13656 13950 13666
rect 14076 13656 14142 13666
rect 14268 13656 14324 13666
rect 14752 13656 14818 13666
rect 14944 13656 15010 13666
rect 15136 13656 15202 13666
rect 15328 13656 15394 13666
rect 15520 13656 15586 13666
rect 15712 13656 15778 13666
rect 15904 13656 15970 13666
rect 16096 13656 16152 13666
rect 16580 13656 16646 13666
rect 16772 13656 16838 13666
rect 16964 13656 17030 13666
rect 17156 13656 17222 13666
rect 17348 13656 17414 13666
rect 17540 13656 17606 13666
rect 17732 13656 17798 13666
rect 17924 13656 17980 13666
rect 18408 13656 18474 13666
rect 18600 13656 18666 13666
rect 18792 13656 18858 13666
rect 18984 13656 19050 13666
rect 19176 13656 19242 13666
rect 19368 13656 19434 13666
rect 19560 13656 19626 13666
rect 19752 13656 19808 13666
rect 20236 13656 20302 13666
rect 20428 13656 20494 13666
rect 20620 13656 20686 13666
rect 20812 13656 20878 13666
rect 21004 13656 21070 13666
rect 21196 13656 21262 13666
rect 21388 13656 21454 13666
rect 21580 13656 21636 13666
rect 32 13318 98 13328
rect 224 13318 290 13328
rect 416 13318 482 13328
rect 608 13318 674 13328
rect 800 13318 866 13328
rect 992 13318 1058 13328
rect 1184 13318 1250 13328
rect 1376 13318 1442 13328
rect 1860 13318 1926 13328
rect 2052 13318 2118 13328
rect 2244 13318 2310 13328
rect 2436 13318 2502 13328
rect 2628 13318 2694 13328
rect 2820 13318 2886 13328
rect 3012 13318 3078 13328
rect 3204 13318 3270 13328
rect 3688 13318 3754 13328
rect 3880 13318 3946 13328
rect 4072 13318 4138 13328
rect 4264 13318 4330 13328
rect 4456 13318 4522 13328
rect 4648 13318 4714 13328
rect 4840 13318 4906 13328
rect 5032 13318 5098 13328
rect 5516 13318 5582 13328
rect 5708 13318 5774 13328
rect 5900 13318 5966 13328
rect 6092 13318 6158 13328
rect 6284 13318 6350 13328
rect 6476 13318 6542 13328
rect 6668 13318 6734 13328
rect 6860 13318 6926 13328
rect 7344 13318 7410 13328
rect 7536 13318 7602 13328
rect 7728 13318 7794 13328
rect 7920 13318 7986 13328
rect 8112 13318 8178 13328
rect 8304 13318 8370 13328
rect 8496 13318 8562 13328
rect 8688 13318 8754 13328
rect 9172 13318 9238 13328
rect 9364 13318 9430 13328
rect 9556 13318 9622 13328
rect 9748 13318 9814 13328
rect 9940 13318 10006 13328
rect 10132 13318 10198 13328
rect 10324 13318 10390 13328
rect 10516 13318 10582 13328
rect 11000 13318 11066 13328
rect 11192 13318 11258 13328
rect 11384 13318 11450 13328
rect 11576 13318 11642 13328
rect 11768 13318 11834 13328
rect 11960 13318 12026 13328
rect 12152 13318 12218 13328
rect 12344 13318 12410 13328
rect 12828 13318 12894 13328
rect 13020 13318 13086 13328
rect 13212 13318 13278 13328
rect 13404 13318 13470 13328
rect 13596 13318 13662 13328
rect 13788 13318 13854 13328
rect 13980 13318 14046 13328
rect 14172 13318 14238 13328
rect 14656 13318 14722 13328
rect 14848 13318 14914 13328
rect 15040 13318 15106 13328
rect 15232 13318 15298 13328
rect 15424 13318 15490 13328
rect 15616 13318 15682 13328
rect 15808 13318 15874 13328
rect 16000 13318 16066 13328
rect 16484 13318 16550 13328
rect 16676 13318 16742 13328
rect 16868 13318 16934 13328
rect 17060 13318 17126 13328
rect 17252 13318 17318 13328
rect 17444 13318 17510 13328
rect 17636 13318 17702 13328
rect 17828 13318 17894 13328
rect 18312 13318 18378 13328
rect 18504 13318 18570 13328
rect 18696 13318 18762 13328
rect 18888 13318 18954 13328
rect 19080 13318 19146 13328
rect 19272 13318 19338 13328
rect 19464 13318 19530 13328
rect 19656 13318 19722 13328
rect 20140 13318 20206 13328
rect 20332 13318 20398 13328
rect 20524 13318 20590 13328
rect 20716 13318 20782 13328
rect 20908 13318 20974 13328
rect 21100 13318 21166 13328
rect 21292 13318 21358 13328
rect 21484 13318 21550 13328
rect 0 13165 32 13318
rect 98 13165 224 13318
rect 290 13165 416 13318
rect 482 13165 608 13318
rect 674 13165 800 13318
rect 866 13165 992 13318
rect 1058 13165 1184 13318
rect 1250 13165 1376 13318
rect 1828 13165 1860 13318
rect 1926 13165 2052 13318
rect 2118 13165 2244 13318
rect 2310 13165 2436 13318
rect 2502 13165 2628 13318
rect 2694 13165 2820 13318
rect 2886 13165 3012 13318
rect 3078 13165 3204 13318
rect 3656 13165 3688 13318
rect 3754 13165 3880 13318
rect 3946 13165 4072 13318
rect 4138 13165 4264 13318
rect 4330 13165 4456 13318
rect 4522 13165 4648 13318
rect 4714 13165 4840 13318
rect 4906 13165 5032 13318
rect 5484 13165 5516 13318
rect 5582 13165 5708 13318
rect 5774 13165 5900 13318
rect 5966 13165 6092 13318
rect 6158 13165 6284 13318
rect 6350 13165 6476 13318
rect 6542 13165 6668 13318
rect 6734 13165 6860 13318
rect 7312 13165 7344 13318
rect 7410 13165 7536 13318
rect 7602 13165 7728 13318
rect 7794 13165 7920 13318
rect 7986 13165 8112 13318
rect 8178 13165 8304 13318
rect 8370 13165 8496 13318
rect 8562 13165 8688 13318
rect 9140 13165 9172 13318
rect 9238 13165 9364 13318
rect 9430 13165 9556 13318
rect 9622 13165 9748 13318
rect 9814 13165 9940 13318
rect 10006 13165 10132 13318
rect 10198 13165 10324 13318
rect 10390 13165 10516 13318
rect 10968 13165 11000 13318
rect 11066 13165 11192 13318
rect 11258 13165 11384 13318
rect 11450 13165 11576 13318
rect 11642 13165 11768 13318
rect 11834 13165 11960 13318
rect 12026 13165 12152 13318
rect 12218 13165 12344 13318
rect 12796 13165 12828 13318
rect 12894 13165 13020 13318
rect 13086 13165 13212 13318
rect 13278 13165 13404 13318
rect 13470 13165 13596 13318
rect 13662 13165 13788 13318
rect 13854 13165 13980 13318
rect 14046 13165 14172 13318
rect 14624 13165 14656 13318
rect 14722 13165 14848 13318
rect 14914 13165 15040 13318
rect 15106 13165 15232 13318
rect 15298 13165 15424 13318
rect 15490 13165 15616 13318
rect 15682 13165 15808 13318
rect 15874 13165 16000 13318
rect 16452 13165 16484 13318
rect 16550 13165 16676 13318
rect 16742 13165 16868 13318
rect 16934 13165 17060 13318
rect 17126 13165 17252 13318
rect 17318 13165 17444 13318
rect 17510 13165 17636 13318
rect 17702 13165 17828 13318
rect 18280 13165 18312 13318
rect 18378 13165 18504 13318
rect 18570 13165 18696 13318
rect 18762 13165 18888 13318
rect 18954 13165 19080 13318
rect 19146 13165 19272 13318
rect 19338 13165 19464 13318
rect 19530 13165 19656 13318
rect 20108 13165 20140 13318
rect 20206 13165 20332 13318
rect 20398 13165 20524 13318
rect 20590 13165 20716 13318
rect 20782 13165 20908 13318
rect 20974 13165 21100 13318
rect 21166 13165 21292 13318
rect 21358 13165 21484 13318
rect 32 13155 98 13165
rect 224 13155 290 13165
rect 416 13155 482 13165
rect 608 13155 674 13165
rect 800 13155 866 13165
rect 992 13155 1058 13165
rect 1184 13155 1250 13165
rect 1376 13155 1442 13165
rect 1860 13155 1926 13165
rect 2052 13155 2118 13165
rect 2244 13155 2310 13165
rect 2436 13155 2502 13165
rect 2628 13155 2694 13165
rect 2820 13155 2886 13165
rect 3012 13155 3078 13165
rect 3204 13155 3270 13165
rect 3688 13155 3754 13165
rect 3880 13155 3946 13165
rect 4072 13155 4138 13165
rect 4264 13155 4330 13165
rect 4456 13155 4522 13165
rect 4648 13155 4714 13165
rect 4840 13155 4906 13165
rect 5032 13155 5098 13165
rect 5516 13155 5582 13165
rect 5708 13155 5774 13165
rect 5900 13155 5966 13165
rect 6092 13155 6158 13165
rect 6284 13155 6350 13165
rect 6476 13155 6542 13165
rect 6668 13155 6734 13165
rect 6860 13155 6926 13165
rect 7344 13155 7410 13165
rect 7536 13155 7602 13165
rect 7728 13155 7794 13165
rect 7920 13155 7986 13165
rect 8112 13155 8178 13165
rect 8304 13155 8370 13165
rect 8496 13155 8562 13165
rect 8688 13155 8754 13165
rect 9172 13155 9238 13165
rect 9364 13155 9430 13165
rect 9556 13155 9622 13165
rect 9748 13155 9814 13165
rect 9940 13155 10006 13165
rect 10132 13155 10198 13165
rect 10324 13155 10390 13165
rect 10516 13155 10582 13165
rect 11000 13155 11066 13165
rect 11192 13155 11258 13165
rect 11384 13155 11450 13165
rect 11576 13155 11642 13165
rect 11768 13155 11834 13165
rect 11960 13155 12026 13165
rect 12152 13155 12218 13165
rect 12344 13155 12410 13165
rect 12828 13155 12894 13165
rect 13020 13155 13086 13165
rect 13212 13155 13278 13165
rect 13404 13155 13470 13165
rect 13596 13155 13662 13165
rect 13788 13155 13854 13165
rect 13980 13155 14046 13165
rect 14172 13155 14238 13165
rect 14656 13155 14722 13165
rect 14848 13155 14914 13165
rect 15040 13155 15106 13165
rect 15232 13155 15298 13165
rect 15424 13155 15490 13165
rect 15616 13155 15682 13165
rect 15808 13155 15874 13165
rect 16000 13155 16066 13165
rect 16484 13155 16550 13165
rect 16676 13155 16742 13165
rect 16868 13155 16934 13165
rect 17060 13155 17126 13165
rect 17252 13155 17318 13165
rect 17444 13155 17510 13165
rect 17636 13155 17702 13165
rect 17828 13155 17894 13165
rect 18312 13155 18378 13165
rect 18504 13155 18570 13165
rect 18696 13155 18762 13165
rect 18888 13155 18954 13165
rect 19080 13155 19146 13165
rect 19272 13155 19338 13165
rect 19464 13155 19530 13165
rect 19656 13155 19722 13165
rect 20140 13155 20206 13165
rect 20332 13155 20398 13165
rect 20524 13155 20590 13165
rect 20716 13155 20782 13165
rect 20908 13155 20974 13165
rect 21100 13155 21166 13165
rect 21292 13155 21358 13165
rect 21484 13155 21550 13165
rect 128 13105 194 13115
rect 320 13105 386 13115
rect 512 13105 578 13115
rect 704 13105 770 13115
rect 896 13105 962 13115
rect 1088 13105 1154 13115
rect 1280 13105 1346 13115
rect 1472 13105 1528 13115
rect 1956 13105 2022 13115
rect 2148 13105 2214 13115
rect 2340 13105 2406 13115
rect 2532 13105 2598 13115
rect 2724 13105 2790 13115
rect 2916 13105 2982 13115
rect 3108 13105 3174 13115
rect 3300 13105 3356 13115
rect 3784 13105 3850 13115
rect 3976 13105 4042 13115
rect 4168 13105 4234 13115
rect 4360 13105 4426 13115
rect 4552 13105 4618 13115
rect 4744 13105 4810 13115
rect 4936 13105 5002 13115
rect 5128 13105 5184 13115
rect 5612 13105 5678 13115
rect 5804 13105 5870 13115
rect 5996 13105 6062 13115
rect 6188 13105 6254 13115
rect 6380 13105 6446 13115
rect 6572 13105 6638 13115
rect 6764 13105 6830 13115
rect 6956 13105 7012 13115
rect 7440 13105 7506 13115
rect 7632 13105 7698 13115
rect 7824 13105 7890 13115
rect 8016 13105 8082 13115
rect 8208 13105 8274 13115
rect 8400 13105 8466 13115
rect 8592 13105 8658 13115
rect 8784 13105 8840 13115
rect 9268 13105 9334 13115
rect 9460 13105 9526 13115
rect 9652 13105 9718 13115
rect 9844 13105 9910 13115
rect 10036 13105 10102 13115
rect 10228 13105 10294 13115
rect 10420 13105 10486 13115
rect 10612 13105 10668 13115
rect 11096 13105 11162 13115
rect 11288 13105 11354 13115
rect 11480 13105 11546 13115
rect 11672 13105 11738 13115
rect 11864 13105 11930 13115
rect 12056 13105 12122 13115
rect 12248 13105 12314 13115
rect 12440 13105 12496 13115
rect 12924 13105 12990 13115
rect 13116 13105 13182 13115
rect 13308 13105 13374 13115
rect 13500 13105 13566 13115
rect 13692 13105 13758 13115
rect 13884 13105 13950 13115
rect 14076 13105 14142 13115
rect 14268 13105 14324 13115
rect 14752 13105 14818 13115
rect 14944 13105 15010 13115
rect 15136 13105 15202 13115
rect 15328 13105 15394 13115
rect 15520 13105 15586 13115
rect 15712 13105 15778 13115
rect 15904 13105 15970 13115
rect 16096 13105 16152 13115
rect 16580 13105 16646 13115
rect 16772 13105 16838 13115
rect 16964 13105 17030 13115
rect 17156 13105 17222 13115
rect 17348 13105 17414 13115
rect 17540 13105 17606 13115
rect 17732 13105 17798 13115
rect 17924 13105 17980 13115
rect 18408 13105 18474 13115
rect 18600 13105 18666 13115
rect 18792 13105 18858 13115
rect 18984 13105 19050 13115
rect 19176 13105 19242 13115
rect 19368 13105 19434 13115
rect 19560 13105 19626 13115
rect 19752 13105 19808 13115
rect 20236 13105 20302 13115
rect 20428 13105 20494 13115
rect 20620 13105 20686 13115
rect 20812 13105 20878 13115
rect 21004 13105 21070 13115
rect 21196 13105 21262 13115
rect 21388 13105 21454 13115
rect 21580 13105 21636 13115
rect 0 12952 128 13105
rect 194 12952 320 13105
rect 386 12952 512 13105
rect 578 12952 704 13105
rect 770 12952 896 13105
rect 962 12952 1088 13105
rect 1154 12952 1280 13105
rect 1346 12952 1472 13105
rect 1528 12952 1708 13105
rect 1828 12952 1956 13105
rect 2022 12952 2148 13105
rect 2214 12952 2340 13105
rect 2406 12952 2532 13105
rect 2598 12952 2724 13105
rect 2790 12952 2916 13105
rect 2982 12952 3108 13105
rect 3174 12952 3300 13105
rect 3356 12952 3536 13105
rect 3656 12952 3784 13105
rect 3850 12952 3976 13105
rect 4042 12952 4168 13105
rect 4234 12952 4360 13105
rect 4426 12952 4552 13105
rect 4618 12952 4744 13105
rect 4810 12952 4936 13105
rect 5002 12952 5128 13105
rect 5184 12952 5364 13105
rect 5484 12952 5612 13105
rect 5678 12952 5804 13105
rect 5870 12952 5996 13105
rect 6062 12952 6188 13105
rect 6254 12952 6380 13105
rect 6446 12952 6572 13105
rect 6638 12952 6764 13105
rect 6830 12952 6956 13105
rect 7012 12952 7192 13105
rect 7312 12952 7440 13105
rect 7506 12952 7632 13105
rect 7698 12952 7824 13105
rect 7890 12952 8016 13105
rect 8082 12952 8208 13105
rect 8274 12952 8400 13105
rect 8466 12952 8592 13105
rect 8658 12952 8784 13105
rect 8840 12952 9020 13105
rect 9140 12952 9268 13105
rect 9334 12952 9460 13105
rect 9526 12952 9652 13105
rect 9718 12952 9844 13105
rect 9910 12952 10036 13105
rect 10102 12952 10228 13105
rect 10294 12952 10420 13105
rect 10486 12952 10612 13105
rect 10668 12952 10848 13105
rect 10968 12952 11096 13105
rect 11162 12952 11288 13105
rect 11354 12952 11480 13105
rect 11546 12952 11672 13105
rect 11738 12952 11864 13105
rect 11930 12952 12056 13105
rect 12122 12952 12248 13105
rect 12314 12952 12440 13105
rect 12496 12952 12676 13105
rect 12796 12952 12924 13105
rect 12990 12952 13116 13105
rect 13182 12952 13308 13105
rect 13374 12952 13500 13105
rect 13566 12952 13692 13105
rect 13758 12952 13884 13105
rect 13950 12952 14076 13105
rect 14142 12952 14268 13105
rect 14324 12952 14504 13105
rect 14624 12952 14752 13105
rect 14818 12952 14944 13105
rect 15010 12952 15136 13105
rect 15202 12952 15328 13105
rect 15394 12952 15520 13105
rect 15586 12952 15712 13105
rect 15778 12952 15904 13105
rect 15970 12952 16096 13105
rect 16152 12952 16332 13105
rect 16452 12952 16580 13105
rect 16646 12952 16772 13105
rect 16838 12952 16964 13105
rect 17030 12952 17156 13105
rect 17222 12952 17348 13105
rect 17414 12952 17540 13105
rect 17606 12952 17732 13105
rect 17798 12952 17924 13105
rect 17980 12952 18160 13105
rect 18280 12952 18408 13105
rect 18474 12952 18600 13105
rect 18666 12952 18792 13105
rect 18858 12952 18984 13105
rect 19050 12952 19176 13105
rect 19242 12952 19368 13105
rect 19434 12952 19560 13105
rect 19626 12952 19752 13105
rect 19808 12952 19988 13105
rect 20108 12952 20236 13105
rect 20302 12952 20428 13105
rect 20494 12952 20620 13105
rect 20686 12952 20812 13105
rect 20878 12952 21004 13105
rect 21070 12952 21196 13105
rect 21262 12952 21388 13105
rect 21454 12952 21580 13105
rect 21636 12952 21816 13105
rect 128 12942 194 12952
rect 320 12942 386 12952
rect 512 12942 578 12952
rect 704 12942 770 12952
rect 896 12942 962 12952
rect 1088 12942 1154 12952
rect 1280 12942 1346 12952
rect 1472 12942 1528 12952
rect 1956 12942 2022 12952
rect 2148 12942 2214 12952
rect 2340 12942 2406 12952
rect 2532 12942 2598 12952
rect 2724 12942 2790 12952
rect 2916 12942 2982 12952
rect 3108 12942 3174 12952
rect 3300 12942 3356 12952
rect 3784 12942 3850 12952
rect 3976 12942 4042 12952
rect 4168 12942 4234 12952
rect 4360 12942 4426 12952
rect 4552 12942 4618 12952
rect 4744 12942 4810 12952
rect 4936 12942 5002 12952
rect 5128 12942 5184 12952
rect 5612 12942 5678 12952
rect 5804 12942 5870 12952
rect 5996 12942 6062 12952
rect 6188 12942 6254 12952
rect 6380 12942 6446 12952
rect 6572 12942 6638 12952
rect 6764 12942 6830 12952
rect 6956 12942 7012 12952
rect 7440 12942 7506 12952
rect 7632 12942 7698 12952
rect 7824 12942 7890 12952
rect 8016 12942 8082 12952
rect 8208 12942 8274 12952
rect 8400 12942 8466 12952
rect 8592 12942 8658 12952
rect 8784 12942 8840 12952
rect 9268 12942 9334 12952
rect 9460 12942 9526 12952
rect 9652 12942 9718 12952
rect 9844 12942 9910 12952
rect 10036 12942 10102 12952
rect 10228 12942 10294 12952
rect 10420 12942 10486 12952
rect 10612 12942 10668 12952
rect 11096 12942 11162 12952
rect 11288 12942 11354 12952
rect 11480 12942 11546 12952
rect 11672 12942 11738 12952
rect 11864 12942 11930 12952
rect 12056 12942 12122 12952
rect 12248 12942 12314 12952
rect 12440 12942 12496 12952
rect 12924 12942 12990 12952
rect 13116 12942 13182 12952
rect 13308 12942 13374 12952
rect 13500 12942 13566 12952
rect 13692 12942 13758 12952
rect 13884 12942 13950 12952
rect 14076 12942 14142 12952
rect 14268 12942 14324 12952
rect 14752 12942 14818 12952
rect 14944 12942 15010 12952
rect 15136 12942 15202 12952
rect 15328 12942 15394 12952
rect 15520 12942 15586 12952
rect 15712 12942 15778 12952
rect 15904 12942 15970 12952
rect 16096 12942 16152 12952
rect 16580 12942 16646 12952
rect 16772 12942 16838 12952
rect 16964 12942 17030 12952
rect 17156 12942 17222 12952
rect 17348 12942 17414 12952
rect 17540 12942 17606 12952
rect 17732 12942 17798 12952
rect 17924 12942 17980 12952
rect 18408 12942 18474 12952
rect 18600 12942 18666 12952
rect 18792 12942 18858 12952
rect 18984 12942 19050 12952
rect 19176 12942 19242 12952
rect 19368 12942 19434 12952
rect 19560 12942 19626 12952
rect 19752 12942 19808 12952
rect 20236 12942 20302 12952
rect 20428 12942 20494 12952
rect 20620 12942 20686 12952
rect 20812 12942 20878 12952
rect 21004 12942 21070 12952
rect 21196 12942 21262 12952
rect 21388 12942 21454 12952
rect 21580 12942 21636 12952
rect 32 12604 98 12614
rect 224 12604 290 12614
rect 416 12604 482 12614
rect 608 12604 674 12614
rect 800 12604 866 12614
rect 992 12604 1058 12614
rect 1184 12604 1250 12614
rect 1376 12604 1442 12614
rect 1860 12604 1926 12614
rect 2052 12604 2118 12614
rect 2244 12604 2310 12614
rect 2436 12604 2502 12614
rect 2628 12604 2694 12614
rect 2820 12604 2886 12614
rect 3012 12604 3078 12614
rect 3204 12604 3270 12614
rect 3688 12604 3754 12614
rect 3880 12604 3946 12614
rect 4072 12604 4138 12614
rect 4264 12604 4330 12614
rect 4456 12604 4522 12614
rect 4648 12604 4714 12614
rect 4840 12604 4906 12614
rect 5032 12604 5098 12614
rect 5516 12604 5582 12614
rect 5708 12604 5774 12614
rect 5900 12604 5966 12614
rect 6092 12604 6158 12614
rect 6284 12604 6350 12614
rect 6476 12604 6542 12614
rect 6668 12604 6734 12614
rect 6860 12604 6926 12614
rect 7344 12604 7410 12614
rect 7536 12604 7602 12614
rect 7728 12604 7794 12614
rect 7920 12604 7986 12614
rect 8112 12604 8178 12614
rect 8304 12604 8370 12614
rect 8496 12604 8562 12614
rect 8688 12604 8754 12614
rect 9172 12604 9238 12614
rect 9364 12604 9430 12614
rect 9556 12604 9622 12614
rect 9748 12604 9814 12614
rect 9940 12604 10006 12614
rect 10132 12604 10198 12614
rect 10324 12604 10390 12614
rect 10516 12604 10582 12614
rect 11000 12604 11066 12614
rect 11192 12604 11258 12614
rect 11384 12604 11450 12614
rect 11576 12604 11642 12614
rect 11768 12604 11834 12614
rect 11960 12604 12026 12614
rect 12152 12604 12218 12614
rect 12344 12604 12410 12614
rect 12828 12604 12894 12614
rect 13020 12604 13086 12614
rect 13212 12604 13278 12614
rect 13404 12604 13470 12614
rect 13596 12604 13662 12614
rect 13788 12604 13854 12614
rect 13980 12604 14046 12614
rect 14172 12604 14238 12614
rect 14656 12604 14722 12614
rect 14848 12604 14914 12614
rect 15040 12604 15106 12614
rect 15232 12604 15298 12614
rect 15424 12604 15490 12614
rect 15616 12604 15682 12614
rect 15808 12604 15874 12614
rect 16000 12604 16066 12614
rect 16484 12604 16550 12614
rect 16676 12604 16742 12614
rect 16868 12604 16934 12614
rect 17060 12604 17126 12614
rect 17252 12604 17318 12614
rect 17444 12604 17510 12614
rect 17636 12604 17702 12614
rect 17828 12604 17894 12614
rect 18312 12604 18378 12614
rect 18504 12604 18570 12614
rect 18696 12604 18762 12614
rect 18888 12604 18954 12614
rect 19080 12604 19146 12614
rect 19272 12604 19338 12614
rect 19464 12604 19530 12614
rect 19656 12604 19722 12614
rect 20140 12604 20206 12614
rect 20332 12604 20398 12614
rect 20524 12604 20590 12614
rect 20716 12604 20782 12614
rect 20908 12604 20974 12614
rect 21100 12604 21166 12614
rect 21292 12604 21358 12614
rect 21484 12604 21550 12614
rect 0 12451 32 12604
rect 98 12451 224 12604
rect 290 12451 416 12604
rect 482 12451 608 12604
rect 674 12451 800 12604
rect 866 12451 992 12604
rect 1058 12451 1184 12604
rect 1250 12451 1376 12604
rect 1828 12451 1860 12604
rect 1926 12451 2052 12604
rect 2118 12451 2244 12604
rect 2310 12451 2436 12604
rect 2502 12451 2628 12604
rect 2694 12451 2820 12604
rect 2886 12451 3012 12604
rect 3078 12451 3204 12604
rect 3656 12451 3688 12604
rect 3754 12451 3880 12604
rect 3946 12451 4072 12604
rect 4138 12451 4264 12604
rect 4330 12451 4456 12604
rect 4522 12451 4648 12604
rect 4714 12451 4840 12604
rect 4906 12451 5032 12604
rect 5484 12451 5516 12604
rect 5582 12451 5708 12604
rect 5774 12451 5900 12604
rect 5966 12451 6092 12604
rect 6158 12451 6284 12604
rect 6350 12451 6476 12604
rect 6542 12451 6668 12604
rect 6734 12451 6860 12604
rect 7312 12451 7344 12604
rect 7410 12451 7536 12604
rect 7602 12451 7728 12604
rect 7794 12451 7920 12604
rect 7986 12451 8112 12604
rect 8178 12451 8304 12604
rect 8370 12451 8496 12604
rect 8562 12451 8688 12604
rect 9140 12451 9172 12604
rect 9238 12451 9364 12604
rect 9430 12451 9556 12604
rect 9622 12451 9748 12604
rect 9814 12451 9940 12604
rect 10006 12451 10132 12604
rect 10198 12451 10324 12604
rect 10390 12451 10516 12604
rect 10968 12451 11000 12604
rect 11066 12451 11192 12604
rect 11258 12451 11384 12604
rect 11450 12451 11576 12604
rect 11642 12451 11768 12604
rect 11834 12451 11960 12604
rect 12026 12451 12152 12604
rect 12218 12451 12344 12604
rect 12796 12451 12828 12604
rect 12894 12451 13020 12604
rect 13086 12451 13212 12604
rect 13278 12451 13404 12604
rect 13470 12451 13596 12604
rect 13662 12451 13788 12604
rect 13854 12451 13980 12604
rect 14046 12451 14172 12604
rect 14624 12451 14656 12604
rect 14722 12451 14848 12604
rect 14914 12451 15040 12604
rect 15106 12451 15232 12604
rect 15298 12451 15424 12604
rect 15490 12451 15616 12604
rect 15682 12451 15808 12604
rect 15874 12451 16000 12604
rect 16452 12451 16484 12604
rect 16550 12451 16676 12604
rect 16742 12451 16868 12604
rect 16934 12451 17060 12604
rect 17126 12451 17252 12604
rect 17318 12451 17444 12604
rect 17510 12451 17636 12604
rect 17702 12451 17828 12604
rect 18280 12451 18312 12604
rect 18378 12451 18504 12604
rect 18570 12451 18696 12604
rect 18762 12451 18888 12604
rect 18954 12451 19080 12604
rect 19146 12451 19272 12604
rect 19338 12451 19464 12604
rect 19530 12451 19656 12604
rect 20108 12451 20140 12604
rect 20206 12451 20332 12604
rect 20398 12451 20524 12604
rect 20590 12451 20716 12604
rect 20782 12451 20908 12604
rect 20974 12451 21100 12604
rect 21166 12451 21292 12604
rect 21358 12451 21484 12604
rect 32 12441 98 12451
rect 224 12441 290 12451
rect 416 12441 482 12451
rect 608 12441 674 12451
rect 800 12441 866 12451
rect 992 12441 1058 12451
rect 1184 12441 1250 12451
rect 1376 12441 1442 12451
rect 1860 12441 1926 12451
rect 2052 12441 2118 12451
rect 2244 12441 2310 12451
rect 2436 12441 2502 12451
rect 2628 12441 2694 12451
rect 2820 12441 2886 12451
rect 3012 12441 3078 12451
rect 3204 12441 3270 12451
rect 3688 12441 3754 12451
rect 3880 12441 3946 12451
rect 4072 12441 4138 12451
rect 4264 12441 4330 12451
rect 4456 12441 4522 12451
rect 4648 12441 4714 12451
rect 4840 12441 4906 12451
rect 5032 12441 5098 12451
rect 5516 12441 5582 12451
rect 5708 12441 5774 12451
rect 5900 12441 5966 12451
rect 6092 12441 6158 12451
rect 6284 12441 6350 12451
rect 6476 12441 6542 12451
rect 6668 12441 6734 12451
rect 6860 12441 6926 12451
rect 7344 12441 7410 12451
rect 7536 12441 7602 12451
rect 7728 12441 7794 12451
rect 7920 12441 7986 12451
rect 8112 12441 8178 12451
rect 8304 12441 8370 12451
rect 8496 12441 8562 12451
rect 8688 12441 8754 12451
rect 9172 12441 9238 12451
rect 9364 12441 9430 12451
rect 9556 12441 9622 12451
rect 9748 12441 9814 12451
rect 9940 12441 10006 12451
rect 10132 12441 10198 12451
rect 10324 12441 10390 12451
rect 10516 12441 10582 12451
rect 11000 12441 11066 12451
rect 11192 12441 11258 12451
rect 11384 12441 11450 12451
rect 11576 12441 11642 12451
rect 11768 12441 11834 12451
rect 11960 12441 12026 12451
rect 12152 12441 12218 12451
rect 12344 12441 12410 12451
rect 12828 12441 12894 12451
rect 13020 12441 13086 12451
rect 13212 12441 13278 12451
rect 13404 12441 13470 12451
rect 13596 12441 13662 12451
rect 13788 12441 13854 12451
rect 13980 12441 14046 12451
rect 14172 12441 14238 12451
rect 14656 12441 14722 12451
rect 14848 12441 14914 12451
rect 15040 12441 15106 12451
rect 15232 12441 15298 12451
rect 15424 12441 15490 12451
rect 15616 12441 15682 12451
rect 15808 12441 15874 12451
rect 16000 12441 16066 12451
rect 16484 12441 16550 12451
rect 16676 12441 16742 12451
rect 16868 12441 16934 12451
rect 17060 12441 17126 12451
rect 17252 12441 17318 12451
rect 17444 12441 17510 12451
rect 17636 12441 17702 12451
rect 17828 12441 17894 12451
rect 18312 12441 18378 12451
rect 18504 12441 18570 12451
rect 18696 12441 18762 12451
rect 18888 12441 18954 12451
rect 19080 12441 19146 12451
rect 19272 12441 19338 12451
rect 19464 12441 19530 12451
rect 19656 12441 19722 12451
rect 20140 12441 20206 12451
rect 20332 12441 20398 12451
rect 20524 12441 20590 12451
rect 20716 12441 20782 12451
rect 20908 12441 20974 12451
rect 21100 12441 21166 12451
rect 21292 12441 21358 12451
rect 21484 12441 21550 12451
rect 128 12391 194 12401
rect 320 12391 386 12401
rect 512 12391 578 12401
rect 704 12391 770 12401
rect 896 12391 962 12401
rect 1088 12391 1154 12401
rect 1280 12391 1346 12401
rect 1472 12391 1528 12401
rect 1956 12391 2022 12401
rect 2148 12391 2214 12401
rect 2340 12391 2406 12401
rect 2532 12391 2598 12401
rect 2724 12391 2790 12401
rect 2916 12391 2982 12401
rect 3108 12391 3174 12401
rect 3300 12391 3356 12401
rect 3784 12391 3850 12401
rect 3976 12391 4042 12401
rect 4168 12391 4234 12401
rect 4360 12391 4426 12401
rect 4552 12391 4618 12401
rect 4744 12391 4810 12401
rect 4936 12391 5002 12401
rect 5128 12391 5184 12401
rect 5612 12391 5678 12401
rect 5804 12391 5870 12401
rect 5996 12391 6062 12401
rect 6188 12391 6254 12401
rect 6380 12391 6446 12401
rect 6572 12391 6638 12401
rect 6764 12391 6830 12401
rect 6956 12391 7012 12401
rect 7440 12391 7506 12401
rect 7632 12391 7698 12401
rect 7824 12391 7890 12401
rect 8016 12391 8082 12401
rect 8208 12391 8274 12401
rect 8400 12391 8466 12401
rect 8592 12391 8658 12401
rect 8784 12391 8840 12401
rect 9268 12391 9334 12401
rect 9460 12391 9526 12401
rect 9652 12391 9718 12401
rect 9844 12391 9910 12401
rect 10036 12391 10102 12401
rect 10228 12391 10294 12401
rect 10420 12391 10486 12401
rect 10612 12391 10668 12401
rect 11096 12391 11162 12401
rect 11288 12391 11354 12401
rect 11480 12391 11546 12401
rect 11672 12391 11738 12401
rect 11864 12391 11930 12401
rect 12056 12391 12122 12401
rect 12248 12391 12314 12401
rect 12440 12391 12496 12401
rect 12924 12391 12990 12401
rect 13116 12391 13182 12401
rect 13308 12391 13374 12401
rect 13500 12391 13566 12401
rect 13692 12391 13758 12401
rect 13884 12391 13950 12401
rect 14076 12391 14142 12401
rect 14268 12391 14324 12401
rect 14752 12391 14818 12401
rect 14944 12391 15010 12401
rect 15136 12391 15202 12401
rect 15328 12391 15394 12401
rect 15520 12391 15586 12401
rect 15712 12391 15778 12401
rect 15904 12391 15970 12401
rect 16096 12391 16152 12401
rect 16580 12391 16646 12401
rect 16772 12391 16838 12401
rect 16964 12391 17030 12401
rect 17156 12391 17222 12401
rect 17348 12391 17414 12401
rect 17540 12391 17606 12401
rect 17732 12391 17798 12401
rect 17924 12391 17980 12401
rect 18408 12391 18474 12401
rect 18600 12391 18666 12401
rect 18792 12391 18858 12401
rect 18984 12391 19050 12401
rect 19176 12391 19242 12401
rect 19368 12391 19434 12401
rect 19560 12391 19626 12401
rect 19752 12391 19808 12401
rect 20236 12391 20302 12401
rect 20428 12391 20494 12401
rect 20620 12391 20686 12401
rect 20812 12391 20878 12401
rect 21004 12391 21070 12401
rect 21196 12391 21262 12401
rect 21388 12391 21454 12401
rect 21580 12391 21636 12401
rect 0 12238 128 12391
rect 194 12238 320 12391
rect 386 12238 512 12391
rect 578 12238 704 12391
rect 770 12238 896 12391
rect 962 12238 1088 12391
rect 1154 12238 1280 12391
rect 1346 12238 1472 12391
rect 1528 12238 1708 12391
rect 1828 12238 1956 12391
rect 2022 12238 2148 12391
rect 2214 12238 2340 12391
rect 2406 12238 2532 12391
rect 2598 12238 2724 12391
rect 2790 12238 2916 12391
rect 2982 12238 3108 12391
rect 3174 12238 3300 12391
rect 3356 12238 3536 12391
rect 3656 12238 3784 12391
rect 3850 12238 3976 12391
rect 4042 12238 4168 12391
rect 4234 12238 4360 12391
rect 4426 12238 4552 12391
rect 4618 12238 4744 12391
rect 4810 12238 4936 12391
rect 5002 12238 5128 12391
rect 5184 12238 5364 12391
rect 5484 12238 5612 12391
rect 5678 12238 5804 12391
rect 5870 12238 5996 12391
rect 6062 12238 6188 12391
rect 6254 12238 6380 12391
rect 6446 12238 6572 12391
rect 6638 12238 6764 12391
rect 6830 12238 6956 12391
rect 7012 12238 7192 12391
rect 7312 12238 7440 12391
rect 7506 12238 7632 12391
rect 7698 12238 7824 12391
rect 7890 12238 8016 12391
rect 8082 12238 8208 12391
rect 8274 12238 8400 12391
rect 8466 12238 8592 12391
rect 8658 12238 8784 12391
rect 8840 12238 9020 12391
rect 9140 12238 9268 12391
rect 9334 12238 9460 12391
rect 9526 12238 9652 12391
rect 9718 12238 9844 12391
rect 9910 12238 10036 12391
rect 10102 12238 10228 12391
rect 10294 12238 10420 12391
rect 10486 12238 10612 12391
rect 10668 12238 10848 12391
rect 10968 12238 11096 12391
rect 11162 12238 11288 12391
rect 11354 12238 11480 12391
rect 11546 12238 11672 12391
rect 11738 12238 11864 12391
rect 11930 12238 12056 12391
rect 12122 12238 12248 12391
rect 12314 12238 12440 12391
rect 12496 12238 12676 12391
rect 12796 12238 12924 12391
rect 12990 12238 13116 12391
rect 13182 12238 13308 12391
rect 13374 12238 13500 12391
rect 13566 12238 13692 12391
rect 13758 12238 13884 12391
rect 13950 12238 14076 12391
rect 14142 12238 14268 12391
rect 14324 12238 14504 12391
rect 14624 12238 14752 12391
rect 14818 12238 14944 12391
rect 15010 12238 15136 12391
rect 15202 12238 15328 12391
rect 15394 12238 15520 12391
rect 15586 12238 15712 12391
rect 15778 12238 15904 12391
rect 15970 12238 16096 12391
rect 16152 12238 16332 12391
rect 16452 12238 16580 12391
rect 16646 12238 16772 12391
rect 16838 12238 16964 12391
rect 17030 12238 17156 12391
rect 17222 12238 17348 12391
rect 17414 12238 17540 12391
rect 17606 12238 17732 12391
rect 17798 12238 17924 12391
rect 17980 12238 18160 12391
rect 18280 12238 18408 12391
rect 18474 12238 18600 12391
rect 18666 12238 18792 12391
rect 18858 12238 18984 12391
rect 19050 12238 19176 12391
rect 19242 12238 19368 12391
rect 19434 12238 19560 12391
rect 19626 12238 19752 12391
rect 19808 12238 19988 12391
rect 20108 12238 20236 12391
rect 20302 12238 20428 12391
rect 20494 12238 20620 12391
rect 20686 12238 20812 12391
rect 20878 12238 21004 12391
rect 21070 12238 21196 12391
rect 21262 12238 21388 12391
rect 21454 12238 21580 12391
rect 21636 12238 21816 12391
rect 128 12228 194 12238
rect 320 12228 386 12238
rect 512 12228 578 12238
rect 704 12228 770 12238
rect 896 12228 962 12238
rect 1088 12228 1154 12238
rect 1280 12228 1346 12238
rect 1472 12228 1528 12238
rect 1956 12228 2022 12238
rect 2148 12228 2214 12238
rect 2340 12228 2406 12238
rect 2532 12228 2598 12238
rect 2724 12228 2790 12238
rect 2916 12228 2982 12238
rect 3108 12228 3174 12238
rect 3300 12228 3356 12238
rect 3784 12228 3850 12238
rect 3976 12228 4042 12238
rect 4168 12228 4234 12238
rect 4360 12228 4426 12238
rect 4552 12228 4618 12238
rect 4744 12228 4810 12238
rect 4936 12228 5002 12238
rect 5128 12228 5184 12238
rect 5612 12228 5678 12238
rect 5804 12228 5870 12238
rect 5996 12228 6062 12238
rect 6188 12228 6254 12238
rect 6380 12228 6446 12238
rect 6572 12228 6638 12238
rect 6764 12228 6830 12238
rect 6956 12228 7012 12238
rect 7440 12228 7506 12238
rect 7632 12228 7698 12238
rect 7824 12228 7890 12238
rect 8016 12228 8082 12238
rect 8208 12228 8274 12238
rect 8400 12228 8466 12238
rect 8592 12228 8658 12238
rect 8784 12228 8840 12238
rect 9268 12228 9334 12238
rect 9460 12228 9526 12238
rect 9652 12228 9718 12238
rect 9844 12228 9910 12238
rect 10036 12228 10102 12238
rect 10228 12228 10294 12238
rect 10420 12228 10486 12238
rect 10612 12228 10668 12238
rect 11096 12228 11162 12238
rect 11288 12228 11354 12238
rect 11480 12228 11546 12238
rect 11672 12228 11738 12238
rect 11864 12228 11930 12238
rect 12056 12228 12122 12238
rect 12248 12228 12314 12238
rect 12440 12228 12496 12238
rect 12924 12228 12990 12238
rect 13116 12228 13182 12238
rect 13308 12228 13374 12238
rect 13500 12228 13566 12238
rect 13692 12228 13758 12238
rect 13884 12228 13950 12238
rect 14076 12228 14142 12238
rect 14268 12228 14324 12238
rect 14752 12228 14818 12238
rect 14944 12228 15010 12238
rect 15136 12228 15202 12238
rect 15328 12228 15394 12238
rect 15520 12228 15586 12238
rect 15712 12228 15778 12238
rect 15904 12228 15970 12238
rect 16096 12228 16152 12238
rect 16580 12228 16646 12238
rect 16772 12228 16838 12238
rect 16964 12228 17030 12238
rect 17156 12228 17222 12238
rect 17348 12228 17414 12238
rect 17540 12228 17606 12238
rect 17732 12228 17798 12238
rect 17924 12228 17980 12238
rect 18408 12228 18474 12238
rect 18600 12228 18666 12238
rect 18792 12228 18858 12238
rect 18984 12228 19050 12238
rect 19176 12228 19242 12238
rect 19368 12228 19434 12238
rect 19560 12228 19626 12238
rect 19752 12228 19808 12238
rect 20236 12228 20302 12238
rect 20428 12228 20494 12238
rect 20620 12228 20686 12238
rect 20812 12228 20878 12238
rect 21004 12228 21070 12238
rect 21196 12228 21262 12238
rect 21388 12228 21454 12238
rect 21580 12228 21636 12238
rect 32 11890 98 11900
rect 224 11890 290 11900
rect 416 11890 482 11900
rect 608 11890 674 11900
rect 800 11890 866 11900
rect 992 11890 1058 11900
rect 1184 11890 1250 11900
rect 1376 11890 1442 11900
rect 1860 11890 1926 11900
rect 2052 11890 2118 11900
rect 2244 11890 2310 11900
rect 2436 11890 2502 11900
rect 2628 11890 2694 11900
rect 2820 11890 2886 11900
rect 3012 11890 3078 11900
rect 3204 11890 3270 11900
rect 3688 11890 3754 11900
rect 3880 11890 3946 11900
rect 4072 11890 4138 11900
rect 4264 11890 4330 11900
rect 4456 11890 4522 11900
rect 4648 11890 4714 11900
rect 4840 11890 4906 11900
rect 5032 11890 5098 11900
rect 5516 11890 5582 11900
rect 5708 11890 5774 11900
rect 5900 11890 5966 11900
rect 6092 11890 6158 11900
rect 6284 11890 6350 11900
rect 6476 11890 6542 11900
rect 6668 11890 6734 11900
rect 6860 11890 6926 11900
rect 7344 11890 7410 11900
rect 7536 11890 7602 11900
rect 7728 11890 7794 11900
rect 7920 11890 7986 11900
rect 8112 11890 8178 11900
rect 8304 11890 8370 11900
rect 8496 11890 8562 11900
rect 8688 11890 8754 11900
rect 9172 11890 9238 11900
rect 9364 11890 9430 11900
rect 9556 11890 9622 11900
rect 9748 11890 9814 11900
rect 9940 11890 10006 11900
rect 10132 11890 10198 11900
rect 10324 11890 10390 11900
rect 10516 11890 10582 11900
rect 11000 11890 11066 11900
rect 11192 11890 11258 11900
rect 11384 11890 11450 11900
rect 11576 11890 11642 11900
rect 11768 11890 11834 11900
rect 11960 11890 12026 11900
rect 12152 11890 12218 11900
rect 12344 11890 12410 11900
rect 12828 11890 12894 11900
rect 13020 11890 13086 11900
rect 13212 11890 13278 11900
rect 13404 11890 13470 11900
rect 13596 11890 13662 11900
rect 13788 11890 13854 11900
rect 13980 11890 14046 11900
rect 14172 11890 14238 11900
rect 14656 11890 14722 11900
rect 14848 11890 14914 11900
rect 15040 11890 15106 11900
rect 15232 11890 15298 11900
rect 15424 11890 15490 11900
rect 15616 11890 15682 11900
rect 15808 11890 15874 11900
rect 16000 11890 16066 11900
rect 16484 11890 16550 11900
rect 16676 11890 16742 11900
rect 16868 11890 16934 11900
rect 17060 11890 17126 11900
rect 17252 11890 17318 11900
rect 17444 11890 17510 11900
rect 17636 11890 17702 11900
rect 17828 11890 17894 11900
rect 18312 11890 18378 11900
rect 18504 11890 18570 11900
rect 18696 11890 18762 11900
rect 18888 11890 18954 11900
rect 19080 11890 19146 11900
rect 19272 11890 19338 11900
rect 19464 11890 19530 11900
rect 19656 11890 19722 11900
rect 20140 11890 20206 11900
rect 20332 11890 20398 11900
rect 20524 11890 20590 11900
rect 20716 11890 20782 11900
rect 20908 11890 20974 11900
rect 21100 11890 21166 11900
rect 21292 11890 21358 11900
rect 21484 11890 21550 11900
rect 0 11737 32 11890
rect 98 11737 224 11890
rect 290 11737 416 11890
rect 482 11737 608 11890
rect 674 11737 800 11890
rect 866 11737 992 11890
rect 1058 11737 1184 11890
rect 1250 11737 1376 11890
rect 1828 11737 1860 11890
rect 1926 11737 2052 11890
rect 2118 11737 2244 11890
rect 2310 11737 2436 11890
rect 2502 11737 2628 11890
rect 2694 11737 2820 11890
rect 2886 11737 3012 11890
rect 3078 11737 3204 11890
rect 3656 11737 3688 11890
rect 3754 11737 3880 11890
rect 3946 11737 4072 11890
rect 4138 11737 4264 11890
rect 4330 11737 4456 11890
rect 4522 11737 4648 11890
rect 4714 11737 4840 11890
rect 4906 11737 5032 11890
rect 5484 11737 5516 11890
rect 5582 11737 5708 11890
rect 5774 11737 5900 11890
rect 5966 11737 6092 11890
rect 6158 11737 6284 11890
rect 6350 11737 6476 11890
rect 6542 11737 6668 11890
rect 6734 11737 6860 11890
rect 7312 11737 7344 11890
rect 7410 11737 7536 11890
rect 7602 11737 7728 11890
rect 7794 11737 7920 11890
rect 7986 11737 8112 11890
rect 8178 11737 8304 11890
rect 8370 11737 8496 11890
rect 8562 11737 8688 11890
rect 9140 11737 9172 11890
rect 9238 11737 9364 11890
rect 9430 11737 9556 11890
rect 9622 11737 9748 11890
rect 9814 11737 9940 11890
rect 10006 11737 10132 11890
rect 10198 11737 10324 11890
rect 10390 11737 10516 11890
rect 10968 11737 11000 11890
rect 11066 11737 11192 11890
rect 11258 11737 11384 11890
rect 11450 11737 11576 11890
rect 11642 11737 11768 11890
rect 11834 11737 11960 11890
rect 12026 11737 12152 11890
rect 12218 11737 12344 11890
rect 12796 11737 12828 11890
rect 12894 11737 13020 11890
rect 13086 11737 13212 11890
rect 13278 11737 13404 11890
rect 13470 11737 13596 11890
rect 13662 11737 13788 11890
rect 13854 11737 13980 11890
rect 14046 11737 14172 11890
rect 14624 11737 14656 11890
rect 14722 11737 14848 11890
rect 14914 11737 15040 11890
rect 15106 11737 15232 11890
rect 15298 11737 15424 11890
rect 15490 11737 15616 11890
rect 15682 11737 15808 11890
rect 15874 11737 16000 11890
rect 16452 11737 16484 11890
rect 16550 11737 16676 11890
rect 16742 11737 16868 11890
rect 16934 11737 17060 11890
rect 17126 11737 17252 11890
rect 17318 11737 17444 11890
rect 17510 11737 17636 11890
rect 17702 11737 17828 11890
rect 18280 11737 18312 11890
rect 18378 11737 18504 11890
rect 18570 11737 18696 11890
rect 18762 11737 18888 11890
rect 18954 11737 19080 11890
rect 19146 11737 19272 11890
rect 19338 11737 19464 11890
rect 19530 11737 19656 11890
rect 20108 11737 20140 11890
rect 20206 11737 20332 11890
rect 20398 11737 20524 11890
rect 20590 11737 20716 11890
rect 20782 11737 20908 11890
rect 20974 11737 21100 11890
rect 21166 11737 21292 11890
rect 21358 11737 21484 11890
rect 32 11727 98 11737
rect 224 11727 290 11737
rect 416 11727 482 11737
rect 608 11727 674 11737
rect 800 11727 866 11737
rect 992 11727 1058 11737
rect 1184 11727 1250 11737
rect 1376 11727 1442 11737
rect 1860 11727 1926 11737
rect 2052 11727 2118 11737
rect 2244 11727 2310 11737
rect 2436 11727 2502 11737
rect 2628 11727 2694 11737
rect 2820 11727 2886 11737
rect 3012 11727 3078 11737
rect 3204 11727 3270 11737
rect 3688 11727 3754 11737
rect 3880 11727 3946 11737
rect 4072 11727 4138 11737
rect 4264 11727 4330 11737
rect 4456 11727 4522 11737
rect 4648 11727 4714 11737
rect 4840 11727 4906 11737
rect 5032 11727 5098 11737
rect 5516 11727 5582 11737
rect 5708 11727 5774 11737
rect 5900 11727 5966 11737
rect 6092 11727 6158 11737
rect 6284 11727 6350 11737
rect 6476 11727 6542 11737
rect 6668 11727 6734 11737
rect 6860 11727 6926 11737
rect 7344 11727 7410 11737
rect 7536 11727 7602 11737
rect 7728 11727 7794 11737
rect 7920 11727 7986 11737
rect 8112 11727 8178 11737
rect 8304 11727 8370 11737
rect 8496 11727 8562 11737
rect 8688 11727 8754 11737
rect 9172 11727 9238 11737
rect 9364 11727 9430 11737
rect 9556 11727 9622 11737
rect 9748 11727 9814 11737
rect 9940 11727 10006 11737
rect 10132 11727 10198 11737
rect 10324 11727 10390 11737
rect 10516 11727 10582 11737
rect 11000 11727 11066 11737
rect 11192 11727 11258 11737
rect 11384 11727 11450 11737
rect 11576 11727 11642 11737
rect 11768 11727 11834 11737
rect 11960 11727 12026 11737
rect 12152 11727 12218 11737
rect 12344 11727 12410 11737
rect 12828 11727 12894 11737
rect 13020 11727 13086 11737
rect 13212 11727 13278 11737
rect 13404 11727 13470 11737
rect 13596 11727 13662 11737
rect 13788 11727 13854 11737
rect 13980 11727 14046 11737
rect 14172 11727 14238 11737
rect 14656 11727 14722 11737
rect 14848 11727 14914 11737
rect 15040 11727 15106 11737
rect 15232 11727 15298 11737
rect 15424 11727 15490 11737
rect 15616 11727 15682 11737
rect 15808 11727 15874 11737
rect 16000 11727 16066 11737
rect 16484 11727 16550 11737
rect 16676 11727 16742 11737
rect 16868 11727 16934 11737
rect 17060 11727 17126 11737
rect 17252 11727 17318 11737
rect 17444 11727 17510 11737
rect 17636 11727 17702 11737
rect 17828 11727 17894 11737
rect 18312 11727 18378 11737
rect 18504 11727 18570 11737
rect 18696 11727 18762 11737
rect 18888 11727 18954 11737
rect 19080 11727 19146 11737
rect 19272 11727 19338 11737
rect 19464 11727 19530 11737
rect 19656 11727 19722 11737
rect 20140 11727 20206 11737
rect 20332 11727 20398 11737
rect 20524 11727 20590 11737
rect 20716 11727 20782 11737
rect 20908 11727 20974 11737
rect 21100 11727 21166 11737
rect 21292 11727 21358 11737
rect 21484 11727 21550 11737
rect 128 11677 194 11687
rect 320 11677 386 11687
rect 512 11677 578 11687
rect 704 11677 770 11687
rect 896 11677 962 11687
rect 1088 11677 1154 11687
rect 1280 11677 1346 11687
rect 1472 11677 1528 11687
rect 1956 11677 2022 11687
rect 2148 11677 2214 11687
rect 2340 11677 2406 11687
rect 2532 11677 2598 11687
rect 2724 11677 2790 11687
rect 2916 11677 2982 11687
rect 3108 11677 3174 11687
rect 3300 11677 3356 11687
rect 3784 11677 3850 11687
rect 3976 11677 4042 11687
rect 4168 11677 4234 11687
rect 4360 11677 4426 11687
rect 4552 11677 4618 11687
rect 4744 11677 4810 11687
rect 4936 11677 5002 11687
rect 5128 11677 5184 11687
rect 5612 11677 5678 11687
rect 5804 11677 5870 11687
rect 5996 11677 6062 11687
rect 6188 11677 6254 11687
rect 6380 11677 6446 11687
rect 6572 11677 6638 11687
rect 6764 11677 6830 11687
rect 6956 11677 7012 11687
rect 7440 11677 7506 11687
rect 7632 11677 7698 11687
rect 7824 11677 7890 11687
rect 8016 11677 8082 11687
rect 8208 11677 8274 11687
rect 8400 11677 8466 11687
rect 8592 11677 8658 11687
rect 8784 11677 8840 11687
rect 9268 11677 9334 11687
rect 9460 11677 9526 11687
rect 9652 11677 9718 11687
rect 9844 11677 9910 11687
rect 10036 11677 10102 11687
rect 10228 11677 10294 11687
rect 10420 11677 10486 11687
rect 10612 11677 10668 11687
rect 11096 11677 11162 11687
rect 11288 11677 11354 11687
rect 11480 11677 11546 11687
rect 11672 11677 11738 11687
rect 11864 11677 11930 11687
rect 12056 11677 12122 11687
rect 12248 11677 12314 11687
rect 12440 11677 12496 11687
rect 12924 11677 12990 11687
rect 13116 11677 13182 11687
rect 13308 11677 13374 11687
rect 13500 11677 13566 11687
rect 13692 11677 13758 11687
rect 13884 11677 13950 11687
rect 14076 11677 14142 11687
rect 14268 11677 14324 11687
rect 14752 11677 14818 11687
rect 14944 11677 15010 11687
rect 15136 11677 15202 11687
rect 15328 11677 15394 11687
rect 15520 11677 15586 11687
rect 15712 11677 15778 11687
rect 15904 11677 15970 11687
rect 16096 11677 16152 11687
rect 16580 11677 16646 11687
rect 16772 11677 16838 11687
rect 16964 11677 17030 11687
rect 17156 11677 17222 11687
rect 17348 11677 17414 11687
rect 17540 11677 17606 11687
rect 17732 11677 17798 11687
rect 17924 11677 17980 11687
rect 18408 11677 18474 11687
rect 18600 11677 18666 11687
rect 18792 11677 18858 11687
rect 18984 11677 19050 11687
rect 19176 11677 19242 11687
rect 19368 11677 19434 11687
rect 19560 11677 19626 11687
rect 19752 11677 19808 11687
rect 20236 11677 20302 11687
rect 20428 11677 20494 11687
rect 20620 11677 20686 11687
rect 20812 11677 20878 11687
rect 21004 11677 21070 11687
rect 21196 11677 21262 11687
rect 21388 11677 21454 11687
rect 21580 11677 21636 11687
rect 0 11524 128 11677
rect 194 11524 320 11677
rect 386 11524 512 11677
rect 578 11524 704 11677
rect 770 11524 896 11677
rect 962 11524 1088 11677
rect 1154 11524 1280 11677
rect 1346 11524 1472 11677
rect 1528 11524 1708 11677
rect 1828 11524 1956 11677
rect 2022 11524 2148 11677
rect 2214 11524 2340 11677
rect 2406 11524 2532 11677
rect 2598 11524 2724 11677
rect 2790 11524 2916 11677
rect 2982 11524 3108 11677
rect 3174 11524 3300 11677
rect 3356 11524 3536 11677
rect 3656 11524 3784 11677
rect 3850 11524 3976 11677
rect 4042 11524 4168 11677
rect 4234 11524 4360 11677
rect 4426 11524 4552 11677
rect 4618 11524 4744 11677
rect 4810 11524 4936 11677
rect 5002 11524 5128 11677
rect 5184 11524 5364 11677
rect 5484 11524 5612 11677
rect 5678 11524 5804 11677
rect 5870 11524 5996 11677
rect 6062 11524 6188 11677
rect 6254 11524 6380 11677
rect 6446 11524 6572 11677
rect 6638 11524 6764 11677
rect 6830 11524 6956 11677
rect 7012 11524 7192 11677
rect 7312 11524 7440 11677
rect 7506 11524 7632 11677
rect 7698 11524 7824 11677
rect 7890 11524 8016 11677
rect 8082 11524 8208 11677
rect 8274 11524 8400 11677
rect 8466 11524 8592 11677
rect 8658 11524 8784 11677
rect 8840 11524 9020 11677
rect 9140 11524 9268 11677
rect 9334 11524 9460 11677
rect 9526 11524 9652 11677
rect 9718 11524 9844 11677
rect 9910 11524 10036 11677
rect 10102 11524 10228 11677
rect 10294 11524 10420 11677
rect 10486 11524 10612 11677
rect 10668 11524 10848 11677
rect 10968 11524 11096 11677
rect 11162 11524 11288 11677
rect 11354 11524 11480 11677
rect 11546 11524 11672 11677
rect 11738 11524 11864 11677
rect 11930 11524 12056 11677
rect 12122 11524 12248 11677
rect 12314 11524 12440 11677
rect 12496 11524 12676 11677
rect 12796 11524 12924 11677
rect 12990 11524 13116 11677
rect 13182 11524 13308 11677
rect 13374 11524 13500 11677
rect 13566 11524 13692 11677
rect 13758 11524 13884 11677
rect 13950 11524 14076 11677
rect 14142 11524 14268 11677
rect 14324 11524 14504 11677
rect 14624 11524 14752 11677
rect 14818 11524 14944 11677
rect 15010 11524 15136 11677
rect 15202 11524 15328 11677
rect 15394 11524 15520 11677
rect 15586 11524 15712 11677
rect 15778 11524 15904 11677
rect 15970 11524 16096 11677
rect 16152 11524 16332 11677
rect 16452 11524 16580 11677
rect 16646 11524 16772 11677
rect 16838 11524 16964 11677
rect 17030 11524 17156 11677
rect 17222 11524 17348 11677
rect 17414 11524 17540 11677
rect 17606 11524 17732 11677
rect 17798 11524 17924 11677
rect 17980 11524 18160 11677
rect 18280 11524 18408 11677
rect 18474 11524 18600 11677
rect 18666 11524 18792 11677
rect 18858 11524 18984 11677
rect 19050 11524 19176 11677
rect 19242 11524 19368 11677
rect 19434 11524 19560 11677
rect 19626 11524 19752 11677
rect 19808 11524 19988 11677
rect 20108 11524 20236 11677
rect 20302 11524 20428 11677
rect 20494 11524 20620 11677
rect 20686 11524 20812 11677
rect 20878 11524 21004 11677
rect 21070 11524 21196 11677
rect 21262 11524 21388 11677
rect 21454 11524 21580 11677
rect 21636 11524 21816 11677
rect 128 11514 194 11524
rect 320 11514 386 11524
rect 512 11514 578 11524
rect 704 11514 770 11524
rect 896 11514 962 11524
rect 1088 11514 1154 11524
rect 1280 11514 1346 11524
rect 1472 11514 1528 11524
rect 1956 11514 2022 11524
rect 2148 11514 2214 11524
rect 2340 11514 2406 11524
rect 2532 11514 2598 11524
rect 2724 11514 2790 11524
rect 2916 11514 2982 11524
rect 3108 11514 3174 11524
rect 3300 11514 3356 11524
rect 3784 11514 3850 11524
rect 3976 11514 4042 11524
rect 4168 11514 4234 11524
rect 4360 11514 4426 11524
rect 4552 11514 4618 11524
rect 4744 11514 4810 11524
rect 4936 11514 5002 11524
rect 5128 11514 5184 11524
rect 5612 11514 5678 11524
rect 5804 11514 5870 11524
rect 5996 11514 6062 11524
rect 6188 11514 6254 11524
rect 6380 11514 6446 11524
rect 6572 11514 6638 11524
rect 6764 11514 6830 11524
rect 6956 11514 7012 11524
rect 7440 11514 7506 11524
rect 7632 11514 7698 11524
rect 7824 11514 7890 11524
rect 8016 11514 8082 11524
rect 8208 11514 8274 11524
rect 8400 11514 8466 11524
rect 8592 11514 8658 11524
rect 8784 11514 8840 11524
rect 9268 11514 9334 11524
rect 9460 11514 9526 11524
rect 9652 11514 9718 11524
rect 9844 11514 9910 11524
rect 10036 11514 10102 11524
rect 10228 11514 10294 11524
rect 10420 11514 10486 11524
rect 10612 11514 10668 11524
rect 11096 11514 11162 11524
rect 11288 11514 11354 11524
rect 11480 11514 11546 11524
rect 11672 11514 11738 11524
rect 11864 11514 11930 11524
rect 12056 11514 12122 11524
rect 12248 11514 12314 11524
rect 12440 11514 12496 11524
rect 12924 11514 12990 11524
rect 13116 11514 13182 11524
rect 13308 11514 13374 11524
rect 13500 11514 13566 11524
rect 13692 11514 13758 11524
rect 13884 11514 13950 11524
rect 14076 11514 14142 11524
rect 14268 11514 14324 11524
rect 14752 11514 14818 11524
rect 14944 11514 15010 11524
rect 15136 11514 15202 11524
rect 15328 11514 15394 11524
rect 15520 11514 15586 11524
rect 15712 11514 15778 11524
rect 15904 11514 15970 11524
rect 16096 11514 16152 11524
rect 16580 11514 16646 11524
rect 16772 11514 16838 11524
rect 16964 11514 17030 11524
rect 17156 11514 17222 11524
rect 17348 11514 17414 11524
rect 17540 11514 17606 11524
rect 17732 11514 17798 11524
rect 17924 11514 17980 11524
rect 18408 11514 18474 11524
rect 18600 11514 18666 11524
rect 18792 11514 18858 11524
rect 18984 11514 19050 11524
rect 19176 11514 19242 11524
rect 19368 11514 19434 11524
rect 19560 11514 19626 11524
rect 19752 11514 19808 11524
rect 20236 11514 20302 11524
rect 20428 11514 20494 11524
rect 20620 11514 20686 11524
rect 20812 11514 20878 11524
rect 21004 11514 21070 11524
rect 21196 11514 21262 11524
rect 21388 11514 21454 11524
rect 21580 11514 21636 11524
rect 32 11176 98 11186
rect 224 11176 290 11186
rect 416 11176 482 11186
rect 608 11176 674 11186
rect 800 11176 866 11186
rect 992 11176 1058 11186
rect 1184 11176 1250 11186
rect 1376 11176 1442 11186
rect 1860 11176 1926 11186
rect 2052 11176 2118 11186
rect 2244 11176 2310 11186
rect 2436 11176 2502 11186
rect 2628 11176 2694 11186
rect 2820 11176 2886 11186
rect 3012 11176 3078 11186
rect 3204 11176 3270 11186
rect 3688 11176 3754 11186
rect 3880 11176 3946 11186
rect 4072 11176 4138 11186
rect 4264 11176 4330 11186
rect 4456 11176 4522 11186
rect 4648 11176 4714 11186
rect 4840 11176 4906 11186
rect 5032 11176 5098 11186
rect 5516 11176 5582 11186
rect 5708 11176 5774 11186
rect 5900 11176 5966 11186
rect 6092 11176 6158 11186
rect 6284 11176 6350 11186
rect 6476 11176 6542 11186
rect 6668 11176 6734 11186
rect 6860 11176 6926 11186
rect 7344 11176 7410 11186
rect 7536 11176 7602 11186
rect 7728 11176 7794 11186
rect 7920 11176 7986 11186
rect 8112 11176 8178 11186
rect 8304 11176 8370 11186
rect 8496 11176 8562 11186
rect 8688 11176 8754 11186
rect 9172 11176 9238 11186
rect 9364 11176 9430 11186
rect 9556 11176 9622 11186
rect 9748 11176 9814 11186
rect 9940 11176 10006 11186
rect 10132 11176 10198 11186
rect 10324 11176 10390 11186
rect 10516 11176 10582 11186
rect 11000 11176 11066 11186
rect 11192 11176 11258 11186
rect 11384 11176 11450 11186
rect 11576 11176 11642 11186
rect 11768 11176 11834 11186
rect 11960 11176 12026 11186
rect 12152 11176 12218 11186
rect 12344 11176 12410 11186
rect 12828 11176 12894 11186
rect 13020 11176 13086 11186
rect 13212 11176 13278 11186
rect 13404 11176 13470 11186
rect 13596 11176 13662 11186
rect 13788 11176 13854 11186
rect 13980 11176 14046 11186
rect 14172 11176 14238 11186
rect 14656 11176 14722 11186
rect 14848 11176 14914 11186
rect 15040 11176 15106 11186
rect 15232 11176 15298 11186
rect 15424 11176 15490 11186
rect 15616 11176 15682 11186
rect 15808 11176 15874 11186
rect 16000 11176 16066 11186
rect 16484 11176 16550 11186
rect 16676 11176 16742 11186
rect 16868 11176 16934 11186
rect 17060 11176 17126 11186
rect 17252 11176 17318 11186
rect 17444 11176 17510 11186
rect 17636 11176 17702 11186
rect 17828 11176 17894 11186
rect 18312 11176 18378 11186
rect 18504 11176 18570 11186
rect 18696 11176 18762 11186
rect 18888 11176 18954 11186
rect 19080 11176 19146 11186
rect 19272 11176 19338 11186
rect 19464 11176 19530 11186
rect 19656 11176 19722 11186
rect 20140 11176 20206 11186
rect 20332 11176 20398 11186
rect 20524 11176 20590 11186
rect 20716 11176 20782 11186
rect 20908 11176 20974 11186
rect 21100 11176 21166 11186
rect 21292 11176 21358 11186
rect 21484 11176 21550 11186
rect 0 11023 32 11176
rect 98 11023 224 11176
rect 290 11023 416 11176
rect 482 11023 608 11176
rect 674 11023 800 11176
rect 866 11023 992 11176
rect 1058 11023 1184 11176
rect 1250 11023 1376 11176
rect 1828 11023 1860 11176
rect 1926 11023 2052 11176
rect 2118 11023 2244 11176
rect 2310 11023 2436 11176
rect 2502 11023 2628 11176
rect 2694 11023 2820 11176
rect 2886 11023 3012 11176
rect 3078 11023 3204 11176
rect 3656 11023 3688 11176
rect 3754 11023 3880 11176
rect 3946 11023 4072 11176
rect 4138 11023 4264 11176
rect 4330 11023 4456 11176
rect 4522 11023 4648 11176
rect 4714 11023 4840 11176
rect 4906 11023 5032 11176
rect 5484 11023 5516 11176
rect 5582 11023 5708 11176
rect 5774 11023 5900 11176
rect 5966 11023 6092 11176
rect 6158 11023 6284 11176
rect 6350 11023 6476 11176
rect 6542 11023 6668 11176
rect 6734 11023 6860 11176
rect 7312 11023 7344 11176
rect 7410 11023 7536 11176
rect 7602 11023 7728 11176
rect 7794 11023 7920 11176
rect 7986 11023 8112 11176
rect 8178 11023 8304 11176
rect 8370 11023 8496 11176
rect 8562 11023 8688 11176
rect 9140 11023 9172 11176
rect 9238 11023 9364 11176
rect 9430 11023 9556 11176
rect 9622 11023 9748 11176
rect 9814 11023 9940 11176
rect 10006 11023 10132 11176
rect 10198 11023 10324 11176
rect 10390 11023 10516 11176
rect 10968 11023 11000 11176
rect 11066 11023 11192 11176
rect 11258 11023 11384 11176
rect 11450 11023 11576 11176
rect 11642 11023 11768 11176
rect 11834 11023 11960 11176
rect 12026 11023 12152 11176
rect 12218 11023 12344 11176
rect 12796 11023 12828 11176
rect 12894 11023 13020 11176
rect 13086 11023 13212 11176
rect 13278 11023 13404 11176
rect 13470 11023 13596 11176
rect 13662 11023 13788 11176
rect 13854 11023 13980 11176
rect 14046 11023 14172 11176
rect 14624 11023 14656 11176
rect 14722 11023 14848 11176
rect 14914 11023 15040 11176
rect 15106 11023 15232 11176
rect 15298 11023 15424 11176
rect 15490 11023 15616 11176
rect 15682 11023 15808 11176
rect 15874 11023 16000 11176
rect 16452 11023 16484 11176
rect 16550 11023 16676 11176
rect 16742 11023 16868 11176
rect 16934 11023 17060 11176
rect 17126 11023 17252 11176
rect 17318 11023 17444 11176
rect 17510 11023 17636 11176
rect 17702 11023 17828 11176
rect 18280 11023 18312 11176
rect 18378 11023 18504 11176
rect 18570 11023 18696 11176
rect 18762 11023 18888 11176
rect 18954 11023 19080 11176
rect 19146 11023 19272 11176
rect 19338 11023 19464 11176
rect 19530 11023 19656 11176
rect 20108 11023 20140 11176
rect 20206 11023 20332 11176
rect 20398 11023 20524 11176
rect 20590 11023 20716 11176
rect 20782 11023 20908 11176
rect 20974 11023 21100 11176
rect 21166 11023 21292 11176
rect 21358 11023 21484 11176
rect 32 11013 98 11023
rect 224 11013 290 11023
rect 416 11013 482 11023
rect 608 11013 674 11023
rect 800 11013 866 11023
rect 992 11013 1058 11023
rect 1184 11013 1250 11023
rect 1376 11013 1442 11023
rect 1860 11013 1926 11023
rect 2052 11013 2118 11023
rect 2244 11013 2310 11023
rect 2436 11013 2502 11023
rect 2628 11013 2694 11023
rect 2820 11013 2886 11023
rect 3012 11013 3078 11023
rect 3204 11013 3270 11023
rect 3688 11013 3754 11023
rect 3880 11013 3946 11023
rect 4072 11013 4138 11023
rect 4264 11013 4330 11023
rect 4456 11013 4522 11023
rect 4648 11013 4714 11023
rect 4840 11013 4906 11023
rect 5032 11013 5098 11023
rect 5516 11013 5582 11023
rect 5708 11013 5774 11023
rect 5900 11013 5966 11023
rect 6092 11013 6158 11023
rect 6284 11013 6350 11023
rect 6476 11013 6542 11023
rect 6668 11013 6734 11023
rect 6860 11013 6926 11023
rect 7344 11013 7410 11023
rect 7536 11013 7602 11023
rect 7728 11013 7794 11023
rect 7920 11013 7986 11023
rect 8112 11013 8178 11023
rect 8304 11013 8370 11023
rect 8496 11013 8562 11023
rect 8688 11013 8754 11023
rect 9172 11013 9238 11023
rect 9364 11013 9430 11023
rect 9556 11013 9622 11023
rect 9748 11013 9814 11023
rect 9940 11013 10006 11023
rect 10132 11013 10198 11023
rect 10324 11013 10390 11023
rect 10516 11013 10582 11023
rect 11000 11013 11066 11023
rect 11192 11013 11258 11023
rect 11384 11013 11450 11023
rect 11576 11013 11642 11023
rect 11768 11013 11834 11023
rect 11960 11013 12026 11023
rect 12152 11013 12218 11023
rect 12344 11013 12410 11023
rect 12828 11013 12894 11023
rect 13020 11013 13086 11023
rect 13212 11013 13278 11023
rect 13404 11013 13470 11023
rect 13596 11013 13662 11023
rect 13788 11013 13854 11023
rect 13980 11013 14046 11023
rect 14172 11013 14238 11023
rect 14656 11013 14722 11023
rect 14848 11013 14914 11023
rect 15040 11013 15106 11023
rect 15232 11013 15298 11023
rect 15424 11013 15490 11023
rect 15616 11013 15682 11023
rect 15808 11013 15874 11023
rect 16000 11013 16066 11023
rect 16484 11013 16550 11023
rect 16676 11013 16742 11023
rect 16868 11013 16934 11023
rect 17060 11013 17126 11023
rect 17252 11013 17318 11023
rect 17444 11013 17510 11023
rect 17636 11013 17702 11023
rect 17828 11013 17894 11023
rect 18312 11013 18378 11023
rect 18504 11013 18570 11023
rect 18696 11013 18762 11023
rect 18888 11013 18954 11023
rect 19080 11013 19146 11023
rect 19272 11013 19338 11023
rect 19464 11013 19530 11023
rect 19656 11013 19722 11023
rect 20140 11013 20206 11023
rect 20332 11013 20398 11023
rect 20524 11013 20590 11023
rect 20716 11013 20782 11023
rect 20908 11013 20974 11023
rect 21100 11013 21166 11023
rect 21292 11013 21358 11023
rect 21484 11013 21550 11023
rect 128 10963 194 10973
rect 320 10963 386 10973
rect 512 10963 578 10973
rect 704 10963 770 10973
rect 896 10963 962 10973
rect 1088 10963 1154 10973
rect 1280 10963 1346 10973
rect 1472 10963 1528 10973
rect 1956 10963 2022 10973
rect 2148 10963 2214 10973
rect 2340 10963 2406 10973
rect 2532 10963 2598 10973
rect 2724 10963 2790 10973
rect 2916 10963 2982 10973
rect 3108 10963 3174 10973
rect 3300 10963 3356 10973
rect 3784 10963 3850 10973
rect 3976 10963 4042 10973
rect 4168 10963 4234 10973
rect 4360 10963 4426 10973
rect 4552 10963 4618 10973
rect 4744 10963 4810 10973
rect 4936 10963 5002 10973
rect 5128 10963 5184 10973
rect 5612 10963 5678 10973
rect 5804 10963 5870 10973
rect 5996 10963 6062 10973
rect 6188 10963 6254 10973
rect 6380 10963 6446 10973
rect 6572 10963 6638 10973
rect 6764 10963 6830 10973
rect 6956 10963 7012 10973
rect 7440 10963 7506 10973
rect 7632 10963 7698 10973
rect 7824 10963 7890 10973
rect 8016 10963 8082 10973
rect 8208 10963 8274 10973
rect 8400 10963 8466 10973
rect 8592 10963 8658 10973
rect 8784 10963 8840 10973
rect 9268 10963 9334 10973
rect 9460 10963 9526 10973
rect 9652 10963 9718 10973
rect 9844 10963 9910 10973
rect 10036 10963 10102 10973
rect 10228 10963 10294 10973
rect 10420 10963 10486 10973
rect 10612 10963 10668 10973
rect 11096 10963 11162 10973
rect 11288 10963 11354 10973
rect 11480 10963 11546 10973
rect 11672 10963 11738 10973
rect 11864 10963 11930 10973
rect 12056 10963 12122 10973
rect 12248 10963 12314 10973
rect 12440 10963 12496 10973
rect 12924 10963 12990 10973
rect 13116 10963 13182 10973
rect 13308 10963 13374 10973
rect 13500 10963 13566 10973
rect 13692 10963 13758 10973
rect 13884 10963 13950 10973
rect 14076 10963 14142 10973
rect 14268 10963 14324 10973
rect 14752 10963 14818 10973
rect 14944 10963 15010 10973
rect 15136 10963 15202 10973
rect 15328 10963 15394 10973
rect 15520 10963 15586 10973
rect 15712 10963 15778 10973
rect 15904 10963 15970 10973
rect 16096 10963 16152 10973
rect 16580 10963 16646 10973
rect 16772 10963 16838 10973
rect 16964 10963 17030 10973
rect 17156 10963 17222 10973
rect 17348 10963 17414 10973
rect 17540 10963 17606 10973
rect 17732 10963 17798 10973
rect 17924 10963 17980 10973
rect 18408 10963 18474 10973
rect 18600 10963 18666 10973
rect 18792 10963 18858 10973
rect 18984 10963 19050 10973
rect 19176 10963 19242 10973
rect 19368 10963 19434 10973
rect 19560 10963 19626 10973
rect 19752 10963 19808 10973
rect 20236 10963 20302 10973
rect 20428 10963 20494 10973
rect 20620 10963 20686 10973
rect 20812 10963 20878 10973
rect 21004 10963 21070 10973
rect 21196 10963 21262 10973
rect 21388 10963 21454 10973
rect 21580 10963 21636 10973
rect 0 10810 128 10963
rect 194 10810 320 10963
rect 386 10810 512 10963
rect 578 10810 704 10963
rect 770 10810 896 10963
rect 962 10810 1088 10963
rect 1154 10810 1280 10963
rect 1346 10810 1472 10963
rect 1528 10810 1708 10963
rect 1828 10810 1956 10963
rect 2022 10810 2148 10963
rect 2214 10810 2340 10963
rect 2406 10810 2532 10963
rect 2598 10810 2724 10963
rect 2790 10810 2916 10963
rect 2982 10810 3108 10963
rect 3174 10810 3300 10963
rect 3356 10810 3536 10963
rect 3656 10810 3784 10963
rect 3850 10810 3976 10963
rect 4042 10810 4168 10963
rect 4234 10810 4360 10963
rect 4426 10810 4552 10963
rect 4618 10810 4744 10963
rect 4810 10810 4936 10963
rect 5002 10810 5128 10963
rect 5184 10810 5364 10963
rect 5484 10810 5612 10963
rect 5678 10810 5804 10963
rect 5870 10810 5996 10963
rect 6062 10810 6188 10963
rect 6254 10810 6380 10963
rect 6446 10810 6572 10963
rect 6638 10810 6764 10963
rect 6830 10810 6956 10963
rect 7012 10810 7192 10963
rect 7312 10810 7440 10963
rect 7506 10810 7632 10963
rect 7698 10810 7824 10963
rect 7890 10810 8016 10963
rect 8082 10810 8208 10963
rect 8274 10810 8400 10963
rect 8466 10810 8592 10963
rect 8658 10810 8784 10963
rect 8840 10810 9020 10963
rect 9140 10810 9268 10963
rect 9334 10810 9460 10963
rect 9526 10810 9652 10963
rect 9718 10810 9844 10963
rect 9910 10810 10036 10963
rect 10102 10810 10228 10963
rect 10294 10810 10420 10963
rect 10486 10810 10612 10963
rect 10668 10810 10848 10963
rect 10968 10810 11096 10963
rect 11162 10810 11288 10963
rect 11354 10810 11480 10963
rect 11546 10810 11672 10963
rect 11738 10810 11864 10963
rect 11930 10810 12056 10963
rect 12122 10810 12248 10963
rect 12314 10810 12440 10963
rect 12496 10810 12676 10963
rect 12796 10810 12924 10963
rect 12990 10810 13116 10963
rect 13182 10810 13308 10963
rect 13374 10810 13500 10963
rect 13566 10810 13692 10963
rect 13758 10810 13884 10963
rect 13950 10810 14076 10963
rect 14142 10810 14268 10963
rect 14324 10810 14504 10963
rect 14624 10810 14752 10963
rect 14818 10810 14944 10963
rect 15010 10810 15136 10963
rect 15202 10810 15328 10963
rect 15394 10810 15520 10963
rect 15586 10810 15712 10963
rect 15778 10810 15904 10963
rect 15970 10810 16096 10963
rect 16152 10810 16332 10963
rect 16452 10810 16580 10963
rect 16646 10810 16772 10963
rect 16838 10810 16964 10963
rect 17030 10810 17156 10963
rect 17222 10810 17348 10963
rect 17414 10810 17540 10963
rect 17606 10810 17732 10963
rect 17798 10810 17924 10963
rect 17980 10810 18160 10963
rect 18280 10810 18408 10963
rect 18474 10810 18600 10963
rect 18666 10810 18792 10963
rect 18858 10810 18984 10963
rect 19050 10810 19176 10963
rect 19242 10810 19368 10963
rect 19434 10810 19560 10963
rect 19626 10810 19752 10963
rect 19808 10810 19988 10963
rect 20108 10810 20236 10963
rect 20302 10810 20428 10963
rect 20494 10810 20620 10963
rect 20686 10810 20812 10963
rect 20878 10810 21004 10963
rect 21070 10810 21196 10963
rect 21262 10810 21388 10963
rect 21454 10810 21580 10963
rect 21636 10810 21816 10963
rect 128 10800 194 10810
rect 320 10800 386 10810
rect 512 10800 578 10810
rect 704 10800 770 10810
rect 896 10800 962 10810
rect 1088 10800 1154 10810
rect 1280 10800 1346 10810
rect 1472 10800 1528 10810
rect 1956 10800 2022 10810
rect 2148 10800 2214 10810
rect 2340 10800 2406 10810
rect 2532 10800 2598 10810
rect 2724 10800 2790 10810
rect 2916 10800 2982 10810
rect 3108 10800 3174 10810
rect 3300 10800 3356 10810
rect 3784 10800 3850 10810
rect 3976 10800 4042 10810
rect 4168 10800 4234 10810
rect 4360 10800 4426 10810
rect 4552 10800 4618 10810
rect 4744 10800 4810 10810
rect 4936 10800 5002 10810
rect 5128 10800 5184 10810
rect 5612 10800 5678 10810
rect 5804 10800 5870 10810
rect 5996 10800 6062 10810
rect 6188 10800 6254 10810
rect 6380 10800 6446 10810
rect 6572 10800 6638 10810
rect 6764 10800 6830 10810
rect 6956 10800 7012 10810
rect 7440 10800 7506 10810
rect 7632 10800 7698 10810
rect 7824 10800 7890 10810
rect 8016 10800 8082 10810
rect 8208 10800 8274 10810
rect 8400 10800 8466 10810
rect 8592 10800 8658 10810
rect 8784 10800 8840 10810
rect 9268 10800 9334 10810
rect 9460 10800 9526 10810
rect 9652 10800 9718 10810
rect 9844 10800 9910 10810
rect 10036 10800 10102 10810
rect 10228 10800 10294 10810
rect 10420 10800 10486 10810
rect 10612 10800 10668 10810
rect 11096 10800 11162 10810
rect 11288 10800 11354 10810
rect 11480 10800 11546 10810
rect 11672 10800 11738 10810
rect 11864 10800 11930 10810
rect 12056 10800 12122 10810
rect 12248 10800 12314 10810
rect 12440 10800 12496 10810
rect 12924 10800 12990 10810
rect 13116 10800 13182 10810
rect 13308 10800 13374 10810
rect 13500 10800 13566 10810
rect 13692 10800 13758 10810
rect 13884 10800 13950 10810
rect 14076 10800 14142 10810
rect 14268 10800 14324 10810
rect 14752 10800 14818 10810
rect 14944 10800 15010 10810
rect 15136 10800 15202 10810
rect 15328 10800 15394 10810
rect 15520 10800 15586 10810
rect 15712 10800 15778 10810
rect 15904 10800 15970 10810
rect 16096 10800 16152 10810
rect 16580 10800 16646 10810
rect 16772 10800 16838 10810
rect 16964 10800 17030 10810
rect 17156 10800 17222 10810
rect 17348 10800 17414 10810
rect 17540 10800 17606 10810
rect 17732 10800 17798 10810
rect 17924 10800 17980 10810
rect 18408 10800 18474 10810
rect 18600 10800 18666 10810
rect 18792 10800 18858 10810
rect 18984 10800 19050 10810
rect 19176 10800 19242 10810
rect 19368 10800 19434 10810
rect 19560 10800 19626 10810
rect 19752 10800 19808 10810
rect 20236 10800 20302 10810
rect 20428 10800 20494 10810
rect 20620 10800 20686 10810
rect 20812 10800 20878 10810
rect 21004 10800 21070 10810
rect 21196 10800 21262 10810
rect 21388 10800 21454 10810
rect 21580 10800 21636 10810
rect 32 10462 98 10472
rect 224 10462 290 10472
rect 416 10462 482 10472
rect 608 10462 674 10472
rect 800 10462 866 10472
rect 992 10462 1058 10472
rect 1184 10462 1250 10472
rect 1376 10462 1442 10472
rect 1860 10462 1926 10472
rect 2052 10462 2118 10472
rect 2244 10462 2310 10472
rect 2436 10462 2502 10472
rect 2628 10462 2694 10472
rect 2820 10462 2886 10472
rect 3012 10462 3078 10472
rect 3204 10462 3270 10472
rect 3688 10462 3754 10472
rect 3880 10462 3946 10472
rect 4072 10462 4138 10472
rect 4264 10462 4330 10472
rect 4456 10462 4522 10472
rect 4648 10462 4714 10472
rect 4840 10462 4906 10472
rect 5032 10462 5098 10472
rect 5516 10462 5582 10472
rect 5708 10462 5774 10472
rect 5900 10462 5966 10472
rect 6092 10462 6158 10472
rect 6284 10462 6350 10472
rect 6476 10462 6542 10472
rect 6668 10462 6734 10472
rect 6860 10462 6926 10472
rect 7344 10462 7410 10472
rect 7536 10462 7602 10472
rect 7728 10462 7794 10472
rect 7920 10462 7986 10472
rect 8112 10462 8178 10472
rect 8304 10462 8370 10472
rect 8496 10462 8562 10472
rect 8688 10462 8754 10472
rect 9172 10462 9238 10472
rect 9364 10462 9430 10472
rect 9556 10462 9622 10472
rect 9748 10462 9814 10472
rect 9940 10462 10006 10472
rect 10132 10462 10198 10472
rect 10324 10462 10390 10472
rect 10516 10462 10582 10472
rect 11000 10462 11066 10472
rect 11192 10462 11258 10472
rect 11384 10462 11450 10472
rect 11576 10462 11642 10472
rect 11768 10462 11834 10472
rect 11960 10462 12026 10472
rect 12152 10462 12218 10472
rect 12344 10462 12410 10472
rect 12828 10462 12894 10472
rect 13020 10462 13086 10472
rect 13212 10462 13278 10472
rect 13404 10462 13470 10472
rect 13596 10462 13662 10472
rect 13788 10462 13854 10472
rect 13980 10462 14046 10472
rect 14172 10462 14238 10472
rect 14656 10462 14722 10472
rect 14848 10462 14914 10472
rect 15040 10462 15106 10472
rect 15232 10462 15298 10472
rect 15424 10462 15490 10472
rect 15616 10462 15682 10472
rect 15808 10462 15874 10472
rect 16000 10462 16066 10472
rect 16484 10462 16550 10472
rect 16676 10462 16742 10472
rect 16868 10462 16934 10472
rect 17060 10462 17126 10472
rect 17252 10462 17318 10472
rect 17444 10462 17510 10472
rect 17636 10462 17702 10472
rect 17828 10462 17894 10472
rect 18312 10462 18378 10472
rect 18504 10462 18570 10472
rect 18696 10462 18762 10472
rect 18888 10462 18954 10472
rect 19080 10462 19146 10472
rect 19272 10462 19338 10472
rect 19464 10462 19530 10472
rect 19656 10462 19722 10472
rect 20140 10462 20206 10472
rect 20332 10462 20398 10472
rect 20524 10462 20590 10472
rect 20716 10462 20782 10472
rect 20908 10462 20974 10472
rect 21100 10462 21166 10472
rect 21292 10462 21358 10472
rect 21484 10462 21550 10472
rect 0 10309 32 10462
rect 98 10309 224 10462
rect 290 10309 416 10462
rect 482 10309 608 10462
rect 674 10309 800 10462
rect 866 10309 992 10462
rect 1058 10309 1184 10462
rect 1250 10309 1376 10462
rect 1828 10309 1860 10462
rect 1926 10309 2052 10462
rect 2118 10309 2244 10462
rect 2310 10309 2436 10462
rect 2502 10309 2628 10462
rect 2694 10309 2820 10462
rect 2886 10309 3012 10462
rect 3078 10309 3204 10462
rect 3656 10309 3688 10462
rect 3754 10309 3880 10462
rect 3946 10309 4072 10462
rect 4138 10309 4264 10462
rect 4330 10309 4456 10462
rect 4522 10309 4648 10462
rect 4714 10309 4840 10462
rect 4906 10309 5032 10462
rect 5484 10309 5516 10462
rect 5582 10309 5708 10462
rect 5774 10309 5900 10462
rect 5966 10309 6092 10462
rect 6158 10309 6284 10462
rect 6350 10309 6476 10462
rect 6542 10309 6668 10462
rect 6734 10309 6860 10462
rect 7312 10309 7344 10462
rect 7410 10309 7536 10462
rect 7602 10309 7728 10462
rect 7794 10309 7920 10462
rect 7986 10309 8112 10462
rect 8178 10309 8304 10462
rect 8370 10309 8496 10462
rect 8562 10309 8688 10462
rect 9140 10309 9172 10462
rect 9238 10309 9364 10462
rect 9430 10309 9556 10462
rect 9622 10309 9748 10462
rect 9814 10309 9940 10462
rect 10006 10309 10132 10462
rect 10198 10309 10324 10462
rect 10390 10309 10516 10462
rect 10968 10309 11000 10462
rect 11066 10309 11192 10462
rect 11258 10309 11384 10462
rect 11450 10309 11576 10462
rect 11642 10309 11768 10462
rect 11834 10309 11960 10462
rect 12026 10309 12152 10462
rect 12218 10309 12344 10462
rect 12796 10309 12828 10462
rect 12894 10309 13020 10462
rect 13086 10309 13212 10462
rect 13278 10309 13404 10462
rect 13470 10309 13596 10462
rect 13662 10309 13788 10462
rect 13854 10309 13980 10462
rect 14046 10309 14172 10462
rect 14624 10309 14656 10462
rect 14722 10309 14848 10462
rect 14914 10309 15040 10462
rect 15106 10309 15232 10462
rect 15298 10309 15424 10462
rect 15490 10309 15616 10462
rect 15682 10309 15808 10462
rect 15874 10309 16000 10462
rect 16452 10309 16484 10462
rect 16550 10309 16676 10462
rect 16742 10309 16868 10462
rect 16934 10309 17060 10462
rect 17126 10309 17252 10462
rect 17318 10309 17444 10462
rect 17510 10309 17636 10462
rect 17702 10309 17828 10462
rect 18280 10309 18312 10462
rect 18378 10309 18504 10462
rect 18570 10309 18696 10462
rect 18762 10309 18888 10462
rect 18954 10309 19080 10462
rect 19146 10309 19272 10462
rect 19338 10309 19464 10462
rect 19530 10309 19656 10462
rect 20108 10309 20140 10462
rect 20206 10309 20332 10462
rect 20398 10309 20524 10462
rect 20590 10309 20716 10462
rect 20782 10309 20908 10462
rect 20974 10309 21100 10462
rect 21166 10309 21292 10462
rect 21358 10309 21484 10462
rect 32 10299 98 10309
rect 224 10299 290 10309
rect 416 10299 482 10309
rect 608 10299 674 10309
rect 800 10299 866 10309
rect 992 10299 1058 10309
rect 1184 10299 1250 10309
rect 1376 10299 1442 10309
rect 1860 10299 1926 10309
rect 2052 10299 2118 10309
rect 2244 10299 2310 10309
rect 2436 10299 2502 10309
rect 2628 10299 2694 10309
rect 2820 10299 2886 10309
rect 3012 10299 3078 10309
rect 3204 10299 3270 10309
rect 3688 10299 3754 10309
rect 3880 10299 3946 10309
rect 4072 10299 4138 10309
rect 4264 10299 4330 10309
rect 4456 10299 4522 10309
rect 4648 10299 4714 10309
rect 4840 10299 4906 10309
rect 5032 10299 5098 10309
rect 5516 10299 5582 10309
rect 5708 10299 5774 10309
rect 5900 10299 5966 10309
rect 6092 10299 6158 10309
rect 6284 10299 6350 10309
rect 6476 10299 6542 10309
rect 6668 10299 6734 10309
rect 6860 10299 6926 10309
rect 7344 10299 7410 10309
rect 7536 10299 7602 10309
rect 7728 10299 7794 10309
rect 7920 10299 7986 10309
rect 8112 10299 8178 10309
rect 8304 10299 8370 10309
rect 8496 10299 8562 10309
rect 8688 10299 8754 10309
rect 9172 10299 9238 10309
rect 9364 10299 9430 10309
rect 9556 10299 9622 10309
rect 9748 10299 9814 10309
rect 9940 10299 10006 10309
rect 10132 10299 10198 10309
rect 10324 10299 10390 10309
rect 10516 10299 10582 10309
rect 11000 10299 11066 10309
rect 11192 10299 11258 10309
rect 11384 10299 11450 10309
rect 11576 10299 11642 10309
rect 11768 10299 11834 10309
rect 11960 10299 12026 10309
rect 12152 10299 12218 10309
rect 12344 10299 12410 10309
rect 12828 10299 12894 10309
rect 13020 10299 13086 10309
rect 13212 10299 13278 10309
rect 13404 10299 13470 10309
rect 13596 10299 13662 10309
rect 13788 10299 13854 10309
rect 13980 10299 14046 10309
rect 14172 10299 14238 10309
rect 14656 10299 14722 10309
rect 14848 10299 14914 10309
rect 15040 10299 15106 10309
rect 15232 10299 15298 10309
rect 15424 10299 15490 10309
rect 15616 10299 15682 10309
rect 15808 10299 15874 10309
rect 16000 10299 16066 10309
rect 16484 10299 16550 10309
rect 16676 10299 16742 10309
rect 16868 10299 16934 10309
rect 17060 10299 17126 10309
rect 17252 10299 17318 10309
rect 17444 10299 17510 10309
rect 17636 10299 17702 10309
rect 17828 10299 17894 10309
rect 18312 10299 18378 10309
rect 18504 10299 18570 10309
rect 18696 10299 18762 10309
rect 18888 10299 18954 10309
rect 19080 10299 19146 10309
rect 19272 10299 19338 10309
rect 19464 10299 19530 10309
rect 19656 10299 19722 10309
rect 20140 10299 20206 10309
rect 20332 10299 20398 10309
rect 20524 10299 20590 10309
rect 20716 10299 20782 10309
rect 20908 10299 20974 10309
rect 21100 10299 21166 10309
rect 21292 10299 21358 10309
rect 21484 10299 21550 10309
rect 128 10249 194 10259
rect 320 10249 386 10259
rect 512 10249 578 10259
rect 704 10249 770 10259
rect 896 10249 962 10259
rect 1088 10249 1154 10259
rect 1280 10249 1346 10259
rect 1472 10249 1528 10259
rect 1956 10249 2022 10259
rect 2148 10249 2214 10259
rect 2340 10249 2406 10259
rect 2532 10249 2598 10259
rect 2724 10249 2790 10259
rect 2916 10249 2982 10259
rect 3108 10249 3174 10259
rect 3300 10249 3356 10259
rect 3784 10249 3850 10259
rect 3976 10249 4042 10259
rect 4168 10249 4234 10259
rect 4360 10249 4426 10259
rect 4552 10249 4618 10259
rect 4744 10249 4810 10259
rect 4936 10249 5002 10259
rect 5128 10249 5184 10259
rect 5612 10249 5678 10259
rect 5804 10249 5870 10259
rect 5996 10249 6062 10259
rect 6188 10249 6254 10259
rect 6380 10249 6446 10259
rect 6572 10249 6638 10259
rect 6764 10249 6830 10259
rect 6956 10249 7012 10259
rect 7440 10249 7506 10259
rect 7632 10249 7698 10259
rect 7824 10249 7890 10259
rect 8016 10249 8082 10259
rect 8208 10249 8274 10259
rect 8400 10249 8466 10259
rect 8592 10249 8658 10259
rect 8784 10249 8840 10259
rect 9268 10249 9334 10259
rect 9460 10249 9526 10259
rect 9652 10249 9718 10259
rect 9844 10249 9910 10259
rect 10036 10249 10102 10259
rect 10228 10249 10294 10259
rect 10420 10249 10486 10259
rect 10612 10249 10668 10259
rect 11096 10249 11162 10259
rect 11288 10249 11354 10259
rect 11480 10249 11546 10259
rect 11672 10249 11738 10259
rect 11864 10249 11930 10259
rect 12056 10249 12122 10259
rect 12248 10249 12314 10259
rect 12440 10249 12496 10259
rect 12924 10249 12990 10259
rect 13116 10249 13182 10259
rect 13308 10249 13374 10259
rect 13500 10249 13566 10259
rect 13692 10249 13758 10259
rect 13884 10249 13950 10259
rect 14076 10249 14142 10259
rect 14268 10249 14324 10259
rect 14752 10249 14818 10259
rect 14944 10249 15010 10259
rect 15136 10249 15202 10259
rect 15328 10249 15394 10259
rect 15520 10249 15586 10259
rect 15712 10249 15778 10259
rect 15904 10249 15970 10259
rect 16096 10249 16152 10259
rect 16580 10249 16646 10259
rect 16772 10249 16838 10259
rect 16964 10249 17030 10259
rect 17156 10249 17222 10259
rect 17348 10249 17414 10259
rect 17540 10249 17606 10259
rect 17732 10249 17798 10259
rect 17924 10249 17980 10259
rect 18408 10249 18474 10259
rect 18600 10249 18666 10259
rect 18792 10249 18858 10259
rect 18984 10249 19050 10259
rect 19176 10249 19242 10259
rect 19368 10249 19434 10259
rect 19560 10249 19626 10259
rect 19752 10249 19808 10259
rect 20236 10249 20302 10259
rect 20428 10249 20494 10259
rect 20620 10249 20686 10259
rect 20812 10249 20878 10259
rect 21004 10249 21070 10259
rect 21196 10249 21262 10259
rect 21388 10249 21454 10259
rect 21580 10249 21636 10259
rect 0 10096 128 10249
rect 194 10096 320 10249
rect 386 10096 512 10249
rect 578 10096 704 10249
rect 770 10096 896 10249
rect 962 10096 1088 10249
rect 1154 10096 1280 10249
rect 1346 10096 1472 10249
rect 1528 10096 1708 10249
rect 1828 10096 1956 10249
rect 2022 10096 2148 10249
rect 2214 10096 2340 10249
rect 2406 10096 2532 10249
rect 2598 10096 2724 10249
rect 2790 10096 2916 10249
rect 2982 10096 3108 10249
rect 3174 10096 3300 10249
rect 3356 10096 3536 10249
rect 3656 10096 3784 10249
rect 3850 10096 3976 10249
rect 4042 10096 4168 10249
rect 4234 10096 4360 10249
rect 4426 10096 4552 10249
rect 4618 10096 4744 10249
rect 4810 10096 4936 10249
rect 5002 10096 5128 10249
rect 5184 10096 5364 10249
rect 5484 10096 5612 10249
rect 5678 10096 5804 10249
rect 5870 10096 5996 10249
rect 6062 10096 6188 10249
rect 6254 10096 6380 10249
rect 6446 10096 6572 10249
rect 6638 10096 6764 10249
rect 6830 10096 6956 10249
rect 7012 10096 7192 10249
rect 7312 10096 7440 10249
rect 7506 10096 7632 10249
rect 7698 10096 7824 10249
rect 7890 10096 8016 10249
rect 8082 10096 8208 10249
rect 8274 10096 8400 10249
rect 8466 10096 8592 10249
rect 8658 10096 8784 10249
rect 8840 10096 9020 10249
rect 9140 10096 9268 10249
rect 9334 10096 9460 10249
rect 9526 10096 9652 10249
rect 9718 10096 9844 10249
rect 9910 10096 10036 10249
rect 10102 10096 10228 10249
rect 10294 10096 10420 10249
rect 10486 10096 10612 10249
rect 10668 10096 10848 10249
rect 10968 10096 11096 10249
rect 11162 10096 11288 10249
rect 11354 10096 11480 10249
rect 11546 10096 11672 10249
rect 11738 10096 11864 10249
rect 11930 10096 12056 10249
rect 12122 10096 12248 10249
rect 12314 10096 12440 10249
rect 12496 10096 12676 10249
rect 12796 10096 12924 10249
rect 12990 10096 13116 10249
rect 13182 10096 13308 10249
rect 13374 10096 13500 10249
rect 13566 10096 13692 10249
rect 13758 10096 13884 10249
rect 13950 10096 14076 10249
rect 14142 10096 14268 10249
rect 14324 10096 14504 10249
rect 14624 10096 14752 10249
rect 14818 10096 14944 10249
rect 15010 10096 15136 10249
rect 15202 10096 15328 10249
rect 15394 10096 15520 10249
rect 15586 10096 15712 10249
rect 15778 10096 15904 10249
rect 15970 10096 16096 10249
rect 16152 10096 16332 10249
rect 16452 10096 16580 10249
rect 16646 10096 16772 10249
rect 16838 10096 16964 10249
rect 17030 10096 17156 10249
rect 17222 10096 17348 10249
rect 17414 10096 17540 10249
rect 17606 10096 17732 10249
rect 17798 10096 17924 10249
rect 17980 10096 18160 10249
rect 18280 10096 18408 10249
rect 18474 10096 18600 10249
rect 18666 10096 18792 10249
rect 18858 10096 18984 10249
rect 19050 10096 19176 10249
rect 19242 10096 19368 10249
rect 19434 10096 19560 10249
rect 19626 10096 19752 10249
rect 19808 10096 19988 10249
rect 20108 10096 20236 10249
rect 20302 10096 20428 10249
rect 20494 10096 20620 10249
rect 20686 10096 20812 10249
rect 20878 10096 21004 10249
rect 21070 10096 21196 10249
rect 21262 10096 21388 10249
rect 21454 10096 21580 10249
rect 21636 10096 21816 10249
rect 128 10086 194 10096
rect 320 10086 386 10096
rect 512 10086 578 10096
rect 704 10086 770 10096
rect 896 10086 962 10096
rect 1088 10086 1154 10096
rect 1280 10086 1346 10096
rect 1472 10086 1528 10096
rect 1956 10086 2022 10096
rect 2148 10086 2214 10096
rect 2340 10086 2406 10096
rect 2532 10086 2598 10096
rect 2724 10086 2790 10096
rect 2916 10086 2982 10096
rect 3108 10086 3174 10096
rect 3300 10086 3356 10096
rect 3784 10086 3850 10096
rect 3976 10086 4042 10096
rect 4168 10086 4234 10096
rect 4360 10086 4426 10096
rect 4552 10086 4618 10096
rect 4744 10086 4810 10096
rect 4936 10086 5002 10096
rect 5128 10086 5184 10096
rect 5612 10086 5678 10096
rect 5804 10086 5870 10096
rect 5996 10086 6062 10096
rect 6188 10086 6254 10096
rect 6380 10086 6446 10096
rect 6572 10086 6638 10096
rect 6764 10086 6830 10096
rect 6956 10086 7012 10096
rect 7440 10086 7506 10096
rect 7632 10086 7698 10096
rect 7824 10086 7890 10096
rect 8016 10086 8082 10096
rect 8208 10086 8274 10096
rect 8400 10086 8466 10096
rect 8592 10086 8658 10096
rect 8784 10086 8840 10096
rect 9268 10086 9334 10096
rect 9460 10086 9526 10096
rect 9652 10086 9718 10096
rect 9844 10086 9910 10096
rect 10036 10086 10102 10096
rect 10228 10086 10294 10096
rect 10420 10086 10486 10096
rect 10612 10086 10668 10096
rect 11096 10086 11162 10096
rect 11288 10086 11354 10096
rect 11480 10086 11546 10096
rect 11672 10086 11738 10096
rect 11864 10086 11930 10096
rect 12056 10086 12122 10096
rect 12248 10086 12314 10096
rect 12440 10086 12496 10096
rect 12924 10086 12990 10096
rect 13116 10086 13182 10096
rect 13308 10086 13374 10096
rect 13500 10086 13566 10096
rect 13692 10086 13758 10096
rect 13884 10086 13950 10096
rect 14076 10086 14142 10096
rect 14268 10086 14324 10096
rect 14752 10086 14818 10096
rect 14944 10086 15010 10096
rect 15136 10086 15202 10096
rect 15328 10086 15394 10096
rect 15520 10086 15586 10096
rect 15712 10086 15778 10096
rect 15904 10086 15970 10096
rect 16096 10086 16152 10096
rect 16580 10086 16646 10096
rect 16772 10086 16838 10096
rect 16964 10086 17030 10096
rect 17156 10086 17222 10096
rect 17348 10086 17414 10096
rect 17540 10086 17606 10096
rect 17732 10086 17798 10096
rect 17924 10086 17980 10096
rect 18408 10086 18474 10096
rect 18600 10086 18666 10096
rect 18792 10086 18858 10096
rect 18984 10086 19050 10096
rect 19176 10086 19242 10096
rect 19368 10086 19434 10096
rect 19560 10086 19626 10096
rect 19752 10086 19808 10096
rect 20236 10086 20302 10096
rect 20428 10086 20494 10096
rect 20620 10086 20686 10096
rect 20812 10086 20878 10096
rect 21004 10086 21070 10096
rect 21196 10086 21262 10096
rect 21388 10086 21454 10096
rect 21580 10086 21636 10096
rect 32 9748 98 9758
rect 224 9748 290 9758
rect 416 9748 482 9758
rect 608 9748 674 9758
rect 800 9748 866 9758
rect 992 9748 1058 9758
rect 1184 9748 1250 9758
rect 1376 9748 1442 9758
rect 1860 9748 1926 9758
rect 2052 9748 2118 9758
rect 2244 9748 2310 9758
rect 2436 9748 2502 9758
rect 2628 9748 2694 9758
rect 2820 9748 2886 9758
rect 3012 9748 3078 9758
rect 3204 9748 3270 9758
rect 3688 9748 3754 9758
rect 3880 9748 3946 9758
rect 4072 9748 4138 9758
rect 4264 9748 4330 9758
rect 4456 9748 4522 9758
rect 4648 9748 4714 9758
rect 4840 9748 4906 9758
rect 5032 9748 5098 9758
rect 5516 9748 5582 9758
rect 5708 9748 5774 9758
rect 5900 9748 5966 9758
rect 6092 9748 6158 9758
rect 6284 9748 6350 9758
rect 6476 9748 6542 9758
rect 6668 9748 6734 9758
rect 6860 9748 6926 9758
rect 7344 9748 7410 9758
rect 7536 9748 7602 9758
rect 7728 9748 7794 9758
rect 7920 9748 7986 9758
rect 8112 9748 8178 9758
rect 8304 9748 8370 9758
rect 8496 9748 8562 9758
rect 8688 9748 8754 9758
rect 9172 9748 9238 9758
rect 9364 9748 9430 9758
rect 9556 9748 9622 9758
rect 9748 9748 9814 9758
rect 9940 9748 10006 9758
rect 10132 9748 10198 9758
rect 10324 9748 10390 9758
rect 10516 9748 10582 9758
rect 11000 9748 11066 9758
rect 11192 9748 11258 9758
rect 11384 9748 11450 9758
rect 11576 9748 11642 9758
rect 11768 9748 11834 9758
rect 11960 9748 12026 9758
rect 12152 9748 12218 9758
rect 12344 9748 12410 9758
rect 12828 9748 12894 9758
rect 13020 9748 13086 9758
rect 13212 9748 13278 9758
rect 13404 9748 13470 9758
rect 13596 9748 13662 9758
rect 13788 9748 13854 9758
rect 13980 9748 14046 9758
rect 14172 9748 14238 9758
rect 14656 9748 14722 9758
rect 14848 9748 14914 9758
rect 15040 9748 15106 9758
rect 15232 9748 15298 9758
rect 15424 9748 15490 9758
rect 15616 9748 15682 9758
rect 15808 9748 15874 9758
rect 16000 9748 16066 9758
rect 16484 9748 16550 9758
rect 16676 9748 16742 9758
rect 16868 9748 16934 9758
rect 17060 9748 17126 9758
rect 17252 9748 17318 9758
rect 17444 9748 17510 9758
rect 17636 9748 17702 9758
rect 17828 9748 17894 9758
rect 18312 9748 18378 9758
rect 18504 9748 18570 9758
rect 18696 9748 18762 9758
rect 18888 9748 18954 9758
rect 19080 9748 19146 9758
rect 19272 9748 19338 9758
rect 19464 9748 19530 9758
rect 19656 9748 19722 9758
rect 20140 9748 20206 9758
rect 20332 9748 20398 9758
rect 20524 9748 20590 9758
rect 20716 9748 20782 9758
rect 20908 9748 20974 9758
rect 21100 9748 21166 9758
rect 21292 9748 21358 9758
rect 21484 9748 21550 9758
rect 0 9595 32 9748
rect 98 9595 224 9748
rect 290 9595 416 9748
rect 482 9595 608 9748
rect 674 9595 800 9748
rect 866 9595 992 9748
rect 1058 9595 1184 9748
rect 1250 9595 1376 9748
rect 1828 9595 1860 9748
rect 1926 9595 2052 9748
rect 2118 9595 2244 9748
rect 2310 9595 2436 9748
rect 2502 9595 2628 9748
rect 2694 9595 2820 9748
rect 2886 9595 3012 9748
rect 3078 9595 3204 9748
rect 3656 9595 3688 9748
rect 3754 9595 3880 9748
rect 3946 9595 4072 9748
rect 4138 9595 4264 9748
rect 4330 9595 4456 9748
rect 4522 9595 4648 9748
rect 4714 9595 4840 9748
rect 4906 9595 5032 9748
rect 5484 9595 5516 9748
rect 5582 9595 5708 9748
rect 5774 9595 5900 9748
rect 5966 9595 6092 9748
rect 6158 9595 6284 9748
rect 6350 9595 6476 9748
rect 6542 9595 6668 9748
rect 6734 9595 6860 9748
rect 7312 9595 7344 9748
rect 7410 9595 7536 9748
rect 7602 9595 7728 9748
rect 7794 9595 7920 9748
rect 7986 9595 8112 9748
rect 8178 9595 8304 9748
rect 8370 9595 8496 9748
rect 8562 9595 8688 9748
rect 9140 9595 9172 9748
rect 9238 9595 9364 9748
rect 9430 9595 9556 9748
rect 9622 9595 9748 9748
rect 9814 9595 9940 9748
rect 10006 9595 10132 9748
rect 10198 9595 10324 9748
rect 10390 9595 10516 9748
rect 10968 9595 11000 9748
rect 11066 9595 11192 9748
rect 11258 9595 11384 9748
rect 11450 9595 11576 9748
rect 11642 9595 11768 9748
rect 11834 9595 11960 9748
rect 12026 9595 12152 9748
rect 12218 9595 12344 9748
rect 12796 9595 12828 9748
rect 12894 9595 13020 9748
rect 13086 9595 13212 9748
rect 13278 9595 13404 9748
rect 13470 9595 13596 9748
rect 13662 9595 13788 9748
rect 13854 9595 13980 9748
rect 14046 9595 14172 9748
rect 14624 9595 14656 9748
rect 14722 9595 14848 9748
rect 14914 9595 15040 9748
rect 15106 9595 15232 9748
rect 15298 9595 15424 9748
rect 15490 9595 15616 9748
rect 15682 9595 15808 9748
rect 15874 9595 16000 9748
rect 16452 9595 16484 9748
rect 16550 9595 16676 9748
rect 16742 9595 16868 9748
rect 16934 9595 17060 9748
rect 17126 9595 17252 9748
rect 17318 9595 17444 9748
rect 17510 9595 17636 9748
rect 17702 9595 17828 9748
rect 18280 9595 18312 9748
rect 18378 9595 18504 9748
rect 18570 9595 18696 9748
rect 18762 9595 18888 9748
rect 18954 9595 19080 9748
rect 19146 9595 19272 9748
rect 19338 9595 19464 9748
rect 19530 9595 19656 9748
rect 20108 9595 20140 9748
rect 20206 9595 20332 9748
rect 20398 9595 20524 9748
rect 20590 9595 20716 9748
rect 20782 9595 20908 9748
rect 20974 9595 21100 9748
rect 21166 9595 21292 9748
rect 21358 9595 21484 9748
rect 32 9585 98 9595
rect 224 9585 290 9595
rect 416 9585 482 9595
rect 608 9585 674 9595
rect 800 9585 866 9595
rect 992 9585 1058 9595
rect 1184 9585 1250 9595
rect 1376 9585 1442 9595
rect 1860 9585 1926 9595
rect 2052 9585 2118 9595
rect 2244 9585 2310 9595
rect 2436 9585 2502 9595
rect 2628 9585 2694 9595
rect 2820 9585 2886 9595
rect 3012 9585 3078 9595
rect 3204 9585 3270 9595
rect 3688 9585 3754 9595
rect 3880 9585 3946 9595
rect 4072 9585 4138 9595
rect 4264 9585 4330 9595
rect 4456 9585 4522 9595
rect 4648 9585 4714 9595
rect 4840 9585 4906 9595
rect 5032 9585 5098 9595
rect 5516 9585 5582 9595
rect 5708 9585 5774 9595
rect 5900 9585 5966 9595
rect 6092 9585 6158 9595
rect 6284 9585 6350 9595
rect 6476 9585 6542 9595
rect 6668 9585 6734 9595
rect 6860 9585 6926 9595
rect 7344 9585 7410 9595
rect 7536 9585 7602 9595
rect 7728 9585 7794 9595
rect 7920 9585 7986 9595
rect 8112 9585 8178 9595
rect 8304 9585 8370 9595
rect 8496 9585 8562 9595
rect 8688 9585 8754 9595
rect 9172 9585 9238 9595
rect 9364 9585 9430 9595
rect 9556 9585 9622 9595
rect 9748 9585 9814 9595
rect 9940 9585 10006 9595
rect 10132 9585 10198 9595
rect 10324 9585 10390 9595
rect 10516 9585 10582 9595
rect 11000 9585 11066 9595
rect 11192 9585 11258 9595
rect 11384 9585 11450 9595
rect 11576 9585 11642 9595
rect 11768 9585 11834 9595
rect 11960 9585 12026 9595
rect 12152 9585 12218 9595
rect 12344 9585 12410 9595
rect 12828 9585 12894 9595
rect 13020 9585 13086 9595
rect 13212 9585 13278 9595
rect 13404 9585 13470 9595
rect 13596 9585 13662 9595
rect 13788 9585 13854 9595
rect 13980 9585 14046 9595
rect 14172 9585 14238 9595
rect 14656 9585 14722 9595
rect 14848 9585 14914 9595
rect 15040 9585 15106 9595
rect 15232 9585 15298 9595
rect 15424 9585 15490 9595
rect 15616 9585 15682 9595
rect 15808 9585 15874 9595
rect 16000 9585 16066 9595
rect 16484 9585 16550 9595
rect 16676 9585 16742 9595
rect 16868 9585 16934 9595
rect 17060 9585 17126 9595
rect 17252 9585 17318 9595
rect 17444 9585 17510 9595
rect 17636 9585 17702 9595
rect 17828 9585 17894 9595
rect 18312 9585 18378 9595
rect 18504 9585 18570 9595
rect 18696 9585 18762 9595
rect 18888 9585 18954 9595
rect 19080 9585 19146 9595
rect 19272 9585 19338 9595
rect 19464 9585 19530 9595
rect 19656 9585 19722 9595
rect 20140 9585 20206 9595
rect 20332 9585 20398 9595
rect 20524 9585 20590 9595
rect 20716 9585 20782 9595
rect 20908 9585 20974 9595
rect 21100 9585 21166 9595
rect 21292 9585 21358 9595
rect 21484 9585 21550 9595
rect 128 9535 194 9545
rect 320 9535 386 9545
rect 512 9535 578 9545
rect 704 9535 770 9545
rect 896 9535 962 9545
rect 1088 9535 1154 9545
rect 1280 9535 1346 9545
rect 1472 9535 1528 9545
rect 1956 9535 2022 9545
rect 2148 9535 2214 9545
rect 2340 9535 2406 9545
rect 2532 9535 2598 9545
rect 2724 9535 2790 9545
rect 2916 9535 2982 9545
rect 3108 9535 3174 9545
rect 3300 9535 3356 9545
rect 3784 9535 3850 9545
rect 3976 9535 4042 9545
rect 4168 9535 4234 9545
rect 4360 9535 4426 9545
rect 4552 9535 4618 9545
rect 4744 9535 4810 9545
rect 4936 9535 5002 9545
rect 5128 9535 5184 9545
rect 5612 9535 5678 9545
rect 5804 9535 5870 9545
rect 5996 9535 6062 9545
rect 6188 9535 6254 9545
rect 6380 9535 6446 9545
rect 6572 9535 6638 9545
rect 6764 9535 6830 9545
rect 6956 9535 7012 9545
rect 7440 9535 7506 9545
rect 7632 9535 7698 9545
rect 7824 9535 7890 9545
rect 8016 9535 8082 9545
rect 8208 9535 8274 9545
rect 8400 9535 8466 9545
rect 8592 9535 8658 9545
rect 8784 9535 8840 9545
rect 9268 9535 9334 9545
rect 9460 9535 9526 9545
rect 9652 9535 9718 9545
rect 9844 9535 9910 9545
rect 10036 9535 10102 9545
rect 10228 9535 10294 9545
rect 10420 9535 10486 9545
rect 10612 9535 10668 9545
rect 11096 9535 11162 9545
rect 11288 9535 11354 9545
rect 11480 9535 11546 9545
rect 11672 9535 11738 9545
rect 11864 9535 11930 9545
rect 12056 9535 12122 9545
rect 12248 9535 12314 9545
rect 12440 9535 12496 9545
rect 12924 9535 12990 9545
rect 13116 9535 13182 9545
rect 13308 9535 13374 9545
rect 13500 9535 13566 9545
rect 13692 9535 13758 9545
rect 13884 9535 13950 9545
rect 14076 9535 14142 9545
rect 14268 9535 14324 9545
rect 14752 9535 14818 9545
rect 14944 9535 15010 9545
rect 15136 9535 15202 9545
rect 15328 9535 15394 9545
rect 15520 9535 15586 9545
rect 15712 9535 15778 9545
rect 15904 9535 15970 9545
rect 16096 9535 16152 9545
rect 16580 9535 16646 9545
rect 16772 9535 16838 9545
rect 16964 9535 17030 9545
rect 17156 9535 17222 9545
rect 17348 9535 17414 9545
rect 17540 9535 17606 9545
rect 17732 9535 17798 9545
rect 17924 9535 17980 9545
rect 18408 9535 18474 9545
rect 18600 9535 18666 9545
rect 18792 9535 18858 9545
rect 18984 9535 19050 9545
rect 19176 9535 19242 9545
rect 19368 9535 19434 9545
rect 19560 9535 19626 9545
rect 19752 9535 19808 9545
rect 20236 9535 20302 9545
rect 20428 9535 20494 9545
rect 20620 9535 20686 9545
rect 20812 9535 20878 9545
rect 21004 9535 21070 9545
rect 21196 9535 21262 9545
rect 21388 9535 21454 9545
rect 21580 9535 21636 9545
rect 0 9382 128 9535
rect 194 9382 320 9535
rect 386 9382 512 9535
rect 578 9382 704 9535
rect 770 9382 896 9535
rect 962 9382 1088 9535
rect 1154 9382 1280 9535
rect 1346 9382 1472 9535
rect 1528 9382 1708 9535
rect 1828 9382 1956 9535
rect 2022 9382 2148 9535
rect 2214 9382 2340 9535
rect 2406 9382 2532 9535
rect 2598 9382 2724 9535
rect 2790 9382 2916 9535
rect 2982 9382 3108 9535
rect 3174 9382 3300 9535
rect 3356 9382 3536 9535
rect 3656 9382 3784 9535
rect 3850 9382 3976 9535
rect 4042 9382 4168 9535
rect 4234 9382 4360 9535
rect 4426 9382 4552 9535
rect 4618 9382 4744 9535
rect 4810 9382 4936 9535
rect 5002 9382 5128 9535
rect 5184 9382 5364 9535
rect 5484 9382 5612 9535
rect 5678 9382 5804 9535
rect 5870 9382 5996 9535
rect 6062 9382 6188 9535
rect 6254 9382 6380 9535
rect 6446 9382 6572 9535
rect 6638 9382 6764 9535
rect 6830 9382 6956 9535
rect 7012 9382 7192 9535
rect 7312 9382 7440 9535
rect 7506 9382 7632 9535
rect 7698 9382 7824 9535
rect 7890 9382 8016 9535
rect 8082 9382 8208 9535
rect 8274 9382 8400 9535
rect 8466 9382 8592 9535
rect 8658 9382 8784 9535
rect 8840 9382 9020 9535
rect 9140 9382 9268 9535
rect 9334 9382 9460 9535
rect 9526 9382 9652 9535
rect 9718 9382 9844 9535
rect 9910 9382 10036 9535
rect 10102 9382 10228 9535
rect 10294 9382 10420 9535
rect 10486 9382 10612 9535
rect 10668 9382 10848 9535
rect 10968 9382 11096 9535
rect 11162 9382 11288 9535
rect 11354 9382 11480 9535
rect 11546 9382 11672 9535
rect 11738 9382 11864 9535
rect 11930 9382 12056 9535
rect 12122 9382 12248 9535
rect 12314 9382 12440 9535
rect 12496 9382 12676 9535
rect 12796 9382 12924 9535
rect 12990 9382 13116 9535
rect 13182 9382 13308 9535
rect 13374 9382 13500 9535
rect 13566 9382 13692 9535
rect 13758 9382 13884 9535
rect 13950 9382 14076 9535
rect 14142 9382 14268 9535
rect 14324 9382 14504 9535
rect 14624 9382 14752 9535
rect 14818 9382 14944 9535
rect 15010 9382 15136 9535
rect 15202 9382 15328 9535
rect 15394 9382 15520 9535
rect 15586 9382 15712 9535
rect 15778 9382 15904 9535
rect 15970 9382 16096 9535
rect 16152 9382 16332 9535
rect 16452 9382 16580 9535
rect 16646 9382 16772 9535
rect 16838 9382 16964 9535
rect 17030 9382 17156 9535
rect 17222 9382 17348 9535
rect 17414 9382 17540 9535
rect 17606 9382 17732 9535
rect 17798 9382 17924 9535
rect 17980 9382 18160 9535
rect 18280 9382 18408 9535
rect 18474 9382 18600 9535
rect 18666 9382 18792 9535
rect 18858 9382 18984 9535
rect 19050 9382 19176 9535
rect 19242 9382 19368 9535
rect 19434 9382 19560 9535
rect 19626 9382 19752 9535
rect 19808 9382 19988 9535
rect 20108 9382 20236 9535
rect 20302 9382 20428 9535
rect 20494 9382 20620 9535
rect 20686 9382 20812 9535
rect 20878 9382 21004 9535
rect 21070 9382 21196 9535
rect 21262 9382 21388 9535
rect 21454 9382 21580 9535
rect 21636 9382 21816 9535
rect 128 9372 194 9382
rect 320 9372 386 9382
rect 512 9372 578 9382
rect 704 9372 770 9382
rect 896 9372 962 9382
rect 1088 9372 1154 9382
rect 1280 9372 1346 9382
rect 1472 9372 1528 9382
rect 1956 9372 2022 9382
rect 2148 9372 2214 9382
rect 2340 9372 2406 9382
rect 2532 9372 2598 9382
rect 2724 9372 2790 9382
rect 2916 9372 2982 9382
rect 3108 9372 3174 9382
rect 3300 9372 3356 9382
rect 3784 9372 3850 9382
rect 3976 9372 4042 9382
rect 4168 9372 4234 9382
rect 4360 9372 4426 9382
rect 4552 9372 4618 9382
rect 4744 9372 4810 9382
rect 4936 9372 5002 9382
rect 5128 9372 5184 9382
rect 5612 9372 5678 9382
rect 5804 9372 5870 9382
rect 5996 9372 6062 9382
rect 6188 9372 6254 9382
rect 6380 9372 6446 9382
rect 6572 9372 6638 9382
rect 6764 9372 6830 9382
rect 6956 9372 7012 9382
rect 7440 9372 7506 9382
rect 7632 9372 7698 9382
rect 7824 9372 7890 9382
rect 8016 9372 8082 9382
rect 8208 9372 8274 9382
rect 8400 9372 8466 9382
rect 8592 9372 8658 9382
rect 8784 9372 8840 9382
rect 9268 9372 9334 9382
rect 9460 9372 9526 9382
rect 9652 9372 9718 9382
rect 9844 9372 9910 9382
rect 10036 9372 10102 9382
rect 10228 9372 10294 9382
rect 10420 9372 10486 9382
rect 10612 9372 10668 9382
rect 11096 9372 11162 9382
rect 11288 9372 11354 9382
rect 11480 9372 11546 9382
rect 11672 9372 11738 9382
rect 11864 9372 11930 9382
rect 12056 9372 12122 9382
rect 12248 9372 12314 9382
rect 12440 9372 12496 9382
rect 12924 9372 12990 9382
rect 13116 9372 13182 9382
rect 13308 9372 13374 9382
rect 13500 9372 13566 9382
rect 13692 9372 13758 9382
rect 13884 9372 13950 9382
rect 14076 9372 14142 9382
rect 14268 9372 14324 9382
rect 14752 9372 14818 9382
rect 14944 9372 15010 9382
rect 15136 9372 15202 9382
rect 15328 9372 15394 9382
rect 15520 9372 15586 9382
rect 15712 9372 15778 9382
rect 15904 9372 15970 9382
rect 16096 9372 16152 9382
rect 16580 9372 16646 9382
rect 16772 9372 16838 9382
rect 16964 9372 17030 9382
rect 17156 9372 17222 9382
rect 17348 9372 17414 9382
rect 17540 9372 17606 9382
rect 17732 9372 17798 9382
rect 17924 9372 17980 9382
rect 18408 9372 18474 9382
rect 18600 9372 18666 9382
rect 18792 9372 18858 9382
rect 18984 9372 19050 9382
rect 19176 9372 19242 9382
rect 19368 9372 19434 9382
rect 19560 9372 19626 9382
rect 19752 9372 19808 9382
rect 20236 9372 20302 9382
rect 20428 9372 20494 9382
rect 20620 9372 20686 9382
rect 20812 9372 20878 9382
rect 21004 9372 21070 9382
rect 21196 9372 21262 9382
rect 21388 9372 21454 9382
rect 21580 9372 21636 9382
rect 32 9034 98 9044
rect 224 9034 290 9044
rect 416 9034 482 9044
rect 608 9034 674 9044
rect 800 9034 866 9044
rect 992 9034 1058 9044
rect 1184 9034 1250 9044
rect 1376 9034 1442 9044
rect 1860 9034 1926 9044
rect 2052 9034 2118 9044
rect 2244 9034 2310 9044
rect 2436 9034 2502 9044
rect 2628 9034 2694 9044
rect 2820 9034 2886 9044
rect 3012 9034 3078 9044
rect 3204 9034 3270 9044
rect 3688 9034 3754 9044
rect 3880 9034 3946 9044
rect 4072 9034 4138 9044
rect 4264 9034 4330 9044
rect 4456 9034 4522 9044
rect 4648 9034 4714 9044
rect 4840 9034 4906 9044
rect 5032 9034 5098 9044
rect 5516 9034 5582 9044
rect 5708 9034 5774 9044
rect 5900 9034 5966 9044
rect 6092 9034 6158 9044
rect 6284 9034 6350 9044
rect 6476 9034 6542 9044
rect 6668 9034 6734 9044
rect 6860 9034 6926 9044
rect 7344 9034 7410 9044
rect 7536 9034 7602 9044
rect 7728 9034 7794 9044
rect 7920 9034 7986 9044
rect 8112 9034 8178 9044
rect 8304 9034 8370 9044
rect 8496 9034 8562 9044
rect 8688 9034 8754 9044
rect 9172 9034 9238 9044
rect 9364 9034 9430 9044
rect 9556 9034 9622 9044
rect 9748 9034 9814 9044
rect 9940 9034 10006 9044
rect 10132 9034 10198 9044
rect 10324 9034 10390 9044
rect 10516 9034 10582 9044
rect 11000 9034 11066 9044
rect 11192 9034 11258 9044
rect 11384 9034 11450 9044
rect 11576 9034 11642 9044
rect 11768 9034 11834 9044
rect 11960 9034 12026 9044
rect 12152 9034 12218 9044
rect 12344 9034 12410 9044
rect 12828 9034 12894 9044
rect 13020 9034 13086 9044
rect 13212 9034 13278 9044
rect 13404 9034 13470 9044
rect 13596 9034 13662 9044
rect 13788 9034 13854 9044
rect 13980 9034 14046 9044
rect 14172 9034 14238 9044
rect 14656 9034 14722 9044
rect 14848 9034 14914 9044
rect 15040 9034 15106 9044
rect 15232 9034 15298 9044
rect 15424 9034 15490 9044
rect 15616 9034 15682 9044
rect 15808 9034 15874 9044
rect 16000 9034 16066 9044
rect 16484 9034 16550 9044
rect 16676 9034 16742 9044
rect 16868 9034 16934 9044
rect 17060 9034 17126 9044
rect 17252 9034 17318 9044
rect 17444 9034 17510 9044
rect 17636 9034 17702 9044
rect 17828 9034 17894 9044
rect 18312 9034 18378 9044
rect 18504 9034 18570 9044
rect 18696 9034 18762 9044
rect 18888 9034 18954 9044
rect 19080 9034 19146 9044
rect 19272 9034 19338 9044
rect 19464 9034 19530 9044
rect 19656 9034 19722 9044
rect 20140 9034 20206 9044
rect 20332 9034 20398 9044
rect 20524 9034 20590 9044
rect 20716 9034 20782 9044
rect 20908 9034 20974 9044
rect 21100 9034 21166 9044
rect 21292 9034 21358 9044
rect 21484 9034 21550 9044
rect 0 8881 32 9034
rect 98 8881 224 9034
rect 290 8881 416 9034
rect 482 8881 608 9034
rect 674 8881 800 9034
rect 866 8881 992 9034
rect 1058 8881 1184 9034
rect 1250 8881 1376 9034
rect 1828 8881 1860 9034
rect 1926 8881 2052 9034
rect 2118 8881 2244 9034
rect 2310 8881 2436 9034
rect 2502 8881 2628 9034
rect 2694 8881 2820 9034
rect 2886 8881 3012 9034
rect 3078 8881 3204 9034
rect 3656 8881 3688 9034
rect 3754 8881 3880 9034
rect 3946 8881 4072 9034
rect 4138 8881 4264 9034
rect 4330 8881 4456 9034
rect 4522 8881 4648 9034
rect 4714 8881 4840 9034
rect 4906 8881 5032 9034
rect 5484 8881 5516 9034
rect 5582 8881 5708 9034
rect 5774 8881 5900 9034
rect 5966 8881 6092 9034
rect 6158 8881 6284 9034
rect 6350 8881 6476 9034
rect 6542 8881 6668 9034
rect 6734 8881 6860 9034
rect 7312 8881 7344 9034
rect 7410 8881 7536 9034
rect 7602 8881 7728 9034
rect 7794 8881 7920 9034
rect 7986 8881 8112 9034
rect 8178 8881 8304 9034
rect 8370 8881 8496 9034
rect 8562 8881 8688 9034
rect 9140 8881 9172 9034
rect 9238 8881 9364 9034
rect 9430 8881 9556 9034
rect 9622 8881 9748 9034
rect 9814 8881 9940 9034
rect 10006 8881 10132 9034
rect 10198 8881 10324 9034
rect 10390 8881 10516 9034
rect 10968 8881 11000 9034
rect 11066 8881 11192 9034
rect 11258 8881 11384 9034
rect 11450 8881 11576 9034
rect 11642 8881 11768 9034
rect 11834 8881 11960 9034
rect 12026 8881 12152 9034
rect 12218 8881 12344 9034
rect 12796 8881 12828 9034
rect 12894 8881 13020 9034
rect 13086 8881 13212 9034
rect 13278 8881 13404 9034
rect 13470 8881 13596 9034
rect 13662 8881 13788 9034
rect 13854 8881 13980 9034
rect 14046 8881 14172 9034
rect 14624 8881 14656 9034
rect 14722 8881 14848 9034
rect 14914 8881 15040 9034
rect 15106 8881 15232 9034
rect 15298 8881 15424 9034
rect 15490 8881 15616 9034
rect 15682 8881 15808 9034
rect 15874 8881 16000 9034
rect 16452 8881 16484 9034
rect 16550 8881 16676 9034
rect 16742 8881 16868 9034
rect 16934 8881 17060 9034
rect 17126 8881 17252 9034
rect 17318 8881 17444 9034
rect 17510 8881 17636 9034
rect 17702 8881 17828 9034
rect 18280 8881 18312 9034
rect 18378 8881 18504 9034
rect 18570 8881 18696 9034
rect 18762 8881 18888 9034
rect 18954 8881 19080 9034
rect 19146 8881 19272 9034
rect 19338 8881 19464 9034
rect 19530 8881 19656 9034
rect 20108 8881 20140 9034
rect 20206 8881 20332 9034
rect 20398 8881 20524 9034
rect 20590 8881 20716 9034
rect 20782 8881 20908 9034
rect 20974 8881 21100 9034
rect 21166 8881 21292 9034
rect 21358 8881 21484 9034
rect 32 8871 98 8881
rect 224 8871 290 8881
rect 416 8871 482 8881
rect 608 8871 674 8881
rect 800 8871 866 8881
rect 992 8871 1058 8881
rect 1184 8871 1250 8881
rect 1376 8871 1442 8881
rect 1860 8871 1926 8881
rect 2052 8871 2118 8881
rect 2244 8871 2310 8881
rect 2436 8871 2502 8881
rect 2628 8871 2694 8881
rect 2820 8871 2886 8881
rect 3012 8871 3078 8881
rect 3204 8871 3270 8881
rect 3688 8871 3754 8881
rect 3880 8871 3946 8881
rect 4072 8871 4138 8881
rect 4264 8871 4330 8881
rect 4456 8871 4522 8881
rect 4648 8871 4714 8881
rect 4840 8871 4906 8881
rect 5032 8871 5098 8881
rect 5516 8871 5582 8881
rect 5708 8871 5774 8881
rect 5900 8871 5966 8881
rect 6092 8871 6158 8881
rect 6284 8871 6350 8881
rect 6476 8871 6542 8881
rect 6668 8871 6734 8881
rect 6860 8871 6926 8881
rect 7344 8871 7410 8881
rect 7536 8871 7602 8881
rect 7728 8871 7794 8881
rect 7920 8871 7986 8881
rect 8112 8871 8178 8881
rect 8304 8871 8370 8881
rect 8496 8871 8562 8881
rect 8688 8871 8754 8881
rect 9172 8871 9238 8881
rect 9364 8871 9430 8881
rect 9556 8871 9622 8881
rect 9748 8871 9814 8881
rect 9940 8871 10006 8881
rect 10132 8871 10198 8881
rect 10324 8871 10390 8881
rect 10516 8871 10582 8881
rect 11000 8871 11066 8881
rect 11192 8871 11258 8881
rect 11384 8871 11450 8881
rect 11576 8871 11642 8881
rect 11768 8871 11834 8881
rect 11960 8871 12026 8881
rect 12152 8871 12218 8881
rect 12344 8871 12410 8881
rect 12828 8871 12894 8881
rect 13020 8871 13086 8881
rect 13212 8871 13278 8881
rect 13404 8871 13470 8881
rect 13596 8871 13662 8881
rect 13788 8871 13854 8881
rect 13980 8871 14046 8881
rect 14172 8871 14238 8881
rect 14656 8871 14722 8881
rect 14848 8871 14914 8881
rect 15040 8871 15106 8881
rect 15232 8871 15298 8881
rect 15424 8871 15490 8881
rect 15616 8871 15682 8881
rect 15808 8871 15874 8881
rect 16000 8871 16066 8881
rect 16484 8871 16550 8881
rect 16676 8871 16742 8881
rect 16868 8871 16934 8881
rect 17060 8871 17126 8881
rect 17252 8871 17318 8881
rect 17444 8871 17510 8881
rect 17636 8871 17702 8881
rect 17828 8871 17894 8881
rect 18312 8871 18378 8881
rect 18504 8871 18570 8881
rect 18696 8871 18762 8881
rect 18888 8871 18954 8881
rect 19080 8871 19146 8881
rect 19272 8871 19338 8881
rect 19464 8871 19530 8881
rect 19656 8871 19722 8881
rect 20140 8871 20206 8881
rect 20332 8871 20398 8881
rect 20524 8871 20590 8881
rect 20716 8871 20782 8881
rect 20908 8871 20974 8881
rect 21100 8871 21166 8881
rect 21292 8871 21358 8881
rect 21484 8871 21550 8881
rect 128 8821 194 8831
rect 320 8821 386 8831
rect 512 8821 578 8831
rect 704 8821 770 8831
rect 896 8821 962 8831
rect 1088 8821 1154 8831
rect 1280 8821 1346 8831
rect 1472 8821 1528 8831
rect 1956 8821 2022 8831
rect 2148 8821 2214 8831
rect 2340 8821 2406 8831
rect 2532 8821 2598 8831
rect 2724 8821 2790 8831
rect 2916 8821 2982 8831
rect 3108 8821 3174 8831
rect 3300 8821 3356 8831
rect 3784 8821 3850 8831
rect 3976 8821 4042 8831
rect 4168 8821 4234 8831
rect 4360 8821 4426 8831
rect 4552 8821 4618 8831
rect 4744 8821 4810 8831
rect 4936 8821 5002 8831
rect 5128 8821 5184 8831
rect 5612 8821 5678 8831
rect 5804 8821 5870 8831
rect 5996 8821 6062 8831
rect 6188 8821 6254 8831
rect 6380 8821 6446 8831
rect 6572 8821 6638 8831
rect 6764 8821 6830 8831
rect 6956 8821 7012 8831
rect 7440 8821 7506 8831
rect 7632 8821 7698 8831
rect 7824 8821 7890 8831
rect 8016 8821 8082 8831
rect 8208 8821 8274 8831
rect 8400 8821 8466 8831
rect 8592 8821 8658 8831
rect 8784 8821 8840 8831
rect 9268 8821 9334 8831
rect 9460 8821 9526 8831
rect 9652 8821 9718 8831
rect 9844 8821 9910 8831
rect 10036 8821 10102 8831
rect 10228 8821 10294 8831
rect 10420 8821 10486 8831
rect 10612 8821 10668 8831
rect 11096 8821 11162 8831
rect 11288 8821 11354 8831
rect 11480 8821 11546 8831
rect 11672 8821 11738 8831
rect 11864 8821 11930 8831
rect 12056 8821 12122 8831
rect 12248 8821 12314 8831
rect 12440 8821 12496 8831
rect 12924 8821 12990 8831
rect 13116 8821 13182 8831
rect 13308 8821 13374 8831
rect 13500 8821 13566 8831
rect 13692 8821 13758 8831
rect 13884 8821 13950 8831
rect 14076 8821 14142 8831
rect 14268 8821 14324 8831
rect 14752 8821 14818 8831
rect 14944 8821 15010 8831
rect 15136 8821 15202 8831
rect 15328 8821 15394 8831
rect 15520 8821 15586 8831
rect 15712 8821 15778 8831
rect 15904 8821 15970 8831
rect 16096 8821 16152 8831
rect 16580 8821 16646 8831
rect 16772 8821 16838 8831
rect 16964 8821 17030 8831
rect 17156 8821 17222 8831
rect 17348 8821 17414 8831
rect 17540 8821 17606 8831
rect 17732 8821 17798 8831
rect 17924 8821 17980 8831
rect 18408 8821 18474 8831
rect 18600 8821 18666 8831
rect 18792 8821 18858 8831
rect 18984 8821 19050 8831
rect 19176 8821 19242 8831
rect 19368 8821 19434 8831
rect 19560 8821 19626 8831
rect 19752 8821 19808 8831
rect 20236 8821 20302 8831
rect 20428 8821 20494 8831
rect 20620 8821 20686 8831
rect 20812 8821 20878 8831
rect 21004 8821 21070 8831
rect 21196 8821 21262 8831
rect 21388 8821 21454 8831
rect 21580 8821 21636 8831
rect 0 8668 128 8821
rect 194 8668 320 8821
rect 386 8668 512 8821
rect 578 8668 704 8821
rect 770 8668 896 8821
rect 962 8668 1088 8821
rect 1154 8668 1280 8821
rect 1346 8668 1472 8821
rect 1528 8668 1708 8821
rect 1828 8668 1956 8821
rect 2022 8668 2148 8821
rect 2214 8668 2340 8821
rect 2406 8668 2532 8821
rect 2598 8668 2724 8821
rect 2790 8668 2916 8821
rect 2982 8668 3108 8821
rect 3174 8668 3300 8821
rect 3356 8668 3536 8821
rect 3656 8668 3784 8821
rect 3850 8668 3976 8821
rect 4042 8668 4168 8821
rect 4234 8668 4360 8821
rect 4426 8668 4552 8821
rect 4618 8668 4744 8821
rect 4810 8668 4936 8821
rect 5002 8668 5128 8821
rect 5184 8668 5364 8821
rect 5484 8668 5612 8821
rect 5678 8668 5804 8821
rect 5870 8668 5996 8821
rect 6062 8668 6188 8821
rect 6254 8668 6380 8821
rect 6446 8668 6572 8821
rect 6638 8668 6764 8821
rect 6830 8668 6956 8821
rect 7012 8668 7192 8821
rect 7312 8668 7440 8821
rect 7506 8668 7632 8821
rect 7698 8668 7824 8821
rect 7890 8668 8016 8821
rect 8082 8668 8208 8821
rect 8274 8668 8400 8821
rect 8466 8668 8592 8821
rect 8658 8668 8784 8821
rect 8840 8668 9020 8821
rect 9140 8668 9268 8821
rect 9334 8668 9460 8821
rect 9526 8668 9652 8821
rect 9718 8668 9844 8821
rect 9910 8668 10036 8821
rect 10102 8668 10228 8821
rect 10294 8668 10420 8821
rect 10486 8668 10612 8821
rect 10668 8668 10848 8821
rect 10968 8668 11096 8821
rect 11162 8668 11288 8821
rect 11354 8668 11480 8821
rect 11546 8668 11672 8821
rect 11738 8668 11864 8821
rect 11930 8668 12056 8821
rect 12122 8668 12248 8821
rect 12314 8668 12440 8821
rect 12496 8668 12676 8821
rect 12796 8668 12924 8821
rect 12990 8668 13116 8821
rect 13182 8668 13308 8821
rect 13374 8668 13500 8821
rect 13566 8668 13692 8821
rect 13758 8668 13884 8821
rect 13950 8668 14076 8821
rect 14142 8668 14268 8821
rect 14324 8668 14504 8821
rect 14624 8668 14752 8821
rect 14818 8668 14944 8821
rect 15010 8668 15136 8821
rect 15202 8668 15328 8821
rect 15394 8668 15520 8821
rect 15586 8668 15712 8821
rect 15778 8668 15904 8821
rect 15970 8668 16096 8821
rect 16152 8668 16332 8821
rect 16452 8668 16580 8821
rect 16646 8668 16772 8821
rect 16838 8668 16964 8821
rect 17030 8668 17156 8821
rect 17222 8668 17348 8821
rect 17414 8668 17540 8821
rect 17606 8668 17732 8821
rect 17798 8668 17924 8821
rect 17980 8668 18160 8821
rect 18280 8668 18408 8821
rect 18474 8668 18600 8821
rect 18666 8668 18792 8821
rect 18858 8668 18984 8821
rect 19050 8668 19176 8821
rect 19242 8668 19368 8821
rect 19434 8668 19560 8821
rect 19626 8668 19752 8821
rect 19808 8668 19988 8821
rect 20108 8668 20236 8821
rect 20302 8668 20428 8821
rect 20494 8668 20620 8821
rect 20686 8668 20812 8821
rect 20878 8668 21004 8821
rect 21070 8668 21196 8821
rect 21262 8668 21388 8821
rect 21454 8668 21580 8821
rect 21636 8668 21816 8821
rect 128 8658 194 8668
rect 320 8658 386 8668
rect 512 8658 578 8668
rect 704 8658 770 8668
rect 896 8658 962 8668
rect 1088 8658 1154 8668
rect 1280 8658 1346 8668
rect 1472 8658 1528 8668
rect 1956 8658 2022 8668
rect 2148 8658 2214 8668
rect 2340 8658 2406 8668
rect 2532 8658 2598 8668
rect 2724 8658 2790 8668
rect 2916 8658 2982 8668
rect 3108 8658 3174 8668
rect 3300 8658 3356 8668
rect 3784 8658 3850 8668
rect 3976 8658 4042 8668
rect 4168 8658 4234 8668
rect 4360 8658 4426 8668
rect 4552 8658 4618 8668
rect 4744 8658 4810 8668
rect 4936 8658 5002 8668
rect 5128 8658 5184 8668
rect 5612 8658 5678 8668
rect 5804 8658 5870 8668
rect 5996 8658 6062 8668
rect 6188 8658 6254 8668
rect 6380 8658 6446 8668
rect 6572 8658 6638 8668
rect 6764 8658 6830 8668
rect 6956 8658 7012 8668
rect 7440 8658 7506 8668
rect 7632 8658 7698 8668
rect 7824 8658 7890 8668
rect 8016 8658 8082 8668
rect 8208 8658 8274 8668
rect 8400 8658 8466 8668
rect 8592 8658 8658 8668
rect 8784 8658 8840 8668
rect 9268 8658 9334 8668
rect 9460 8658 9526 8668
rect 9652 8658 9718 8668
rect 9844 8658 9910 8668
rect 10036 8658 10102 8668
rect 10228 8658 10294 8668
rect 10420 8658 10486 8668
rect 10612 8658 10668 8668
rect 11096 8658 11162 8668
rect 11288 8658 11354 8668
rect 11480 8658 11546 8668
rect 11672 8658 11738 8668
rect 11864 8658 11930 8668
rect 12056 8658 12122 8668
rect 12248 8658 12314 8668
rect 12440 8658 12496 8668
rect 12924 8658 12990 8668
rect 13116 8658 13182 8668
rect 13308 8658 13374 8668
rect 13500 8658 13566 8668
rect 13692 8658 13758 8668
rect 13884 8658 13950 8668
rect 14076 8658 14142 8668
rect 14268 8658 14324 8668
rect 14752 8658 14818 8668
rect 14944 8658 15010 8668
rect 15136 8658 15202 8668
rect 15328 8658 15394 8668
rect 15520 8658 15586 8668
rect 15712 8658 15778 8668
rect 15904 8658 15970 8668
rect 16096 8658 16152 8668
rect 16580 8658 16646 8668
rect 16772 8658 16838 8668
rect 16964 8658 17030 8668
rect 17156 8658 17222 8668
rect 17348 8658 17414 8668
rect 17540 8658 17606 8668
rect 17732 8658 17798 8668
rect 17924 8658 17980 8668
rect 18408 8658 18474 8668
rect 18600 8658 18666 8668
rect 18792 8658 18858 8668
rect 18984 8658 19050 8668
rect 19176 8658 19242 8668
rect 19368 8658 19434 8668
rect 19560 8658 19626 8668
rect 19752 8658 19808 8668
rect 20236 8658 20302 8668
rect 20428 8658 20494 8668
rect 20620 8658 20686 8668
rect 20812 8658 20878 8668
rect 21004 8658 21070 8668
rect 21196 8658 21262 8668
rect 21388 8658 21454 8668
rect 21580 8658 21636 8668
rect 32 8320 98 8330
rect 224 8320 290 8330
rect 416 8320 482 8330
rect 608 8320 674 8330
rect 800 8320 866 8330
rect 992 8320 1058 8330
rect 1184 8320 1250 8330
rect 1376 8320 1442 8330
rect 1860 8320 1926 8330
rect 2052 8320 2118 8330
rect 2244 8320 2310 8330
rect 2436 8320 2502 8330
rect 2628 8320 2694 8330
rect 2820 8320 2886 8330
rect 3012 8320 3078 8330
rect 3204 8320 3270 8330
rect 3688 8320 3754 8330
rect 3880 8320 3946 8330
rect 4072 8320 4138 8330
rect 4264 8320 4330 8330
rect 4456 8320 4522 8330
rect 4648 8320 4714 8330
rect 4840 8320 4906 8330
rect 5032 8320 5098 8330
rect 5516 8320 5582 8330
rect 5708 8320 5774 8330
rect 5900 8320 5966 8330
rect 6092 8320 6158 8330
rect 6284 8320 6350 8330
rect 6476 8320 6542 8330
rect 6668 8320 6734 8330
rect 6860 8320 6926 8330
rect 7344 8320 7410 8330
rect 7536 8320 7602 8330
rect 7728 8320 7794 8330
rect 7920 8320 7986 8330
rect 8112 8320 8178 8330
rect 8304 8320 8370 8330
rect 8496 8320 8562 8330
rect 8688 8320 8754 8330
rect 9172 8320 9238 8330
rect 9364 8320 9430 8330
rect 9556 8320 9622 8330
rect 9748 8320 9814 8330
rect 9940 8320 10006 8330
rect 10132 8320 10198 8330
rect 10324 8320 10390 8330
rect 10516 8320 10582 8330
rect 11000 8320 11066 8330
rect 11192 8320 11258 8330
rect 11384 8320 11450 8330
rect 11576 8320 11642 8330
rect 11768 8320 11834 8330
rect 11960 8320 12026 8330
rect 12152 8320 12218 8330
rect 12344 8320 12410 8330
rect 12828 8320 12894 8330
rect 13020 8320 13086 8330
rect 13212 8320 13278 8330
rect 13404 8320 13470 8330
rect 13596 8320 13662 8330
rect 13788 8320 13854 8330
rect 13980 8320 14046 8330
rect 14172 8320 14238 8330
rect 14656 8320 14722 8330
rect 14848 8320 14914 8330
rect 15040 8320 15106 8330
rect 15232 8320 15298 8330
rect 15424 8320 15490 8330
rect 15616 8320 15682 8330
rect 15808 8320 15874 8330
rect 16000 8320 16066 8330
rect 16484 8320 16550 8330
rect 16676 8320 16742 8330
rect 16868 8320 16934 8330
rect 17060 8320 17126 8330
rect 17252 8320 17318 8330
rect 17444 8320 17510 8330
rect 17636 8320 17702 8330
rect 17828 8320 17894 8330
rect 18312 8320 18378 8330
rect 18504 8320 18570 8330
rect 18696 8320 18762 8330
rect 18888 8320 18954 8330
rect 19080 8320 19146 8330
rect 19272 8320 19338 8330
rect 19464 8320 19530 8330
rect 19656 8320 19722 8330
rect 20140 8320 20206 8330
rect 20332 8320 20398 8330
rect 20524 8320 20590 8330
rect 20716 8320 20782 8330
rect 20908 8320 20974 8330
rect 21100 8320 21166 8330
rect 21292 8320 21358 8330
rect 21484 8320 21550 8330
rect 0 8167 32 8320
rect 98 8167 224 8320
rect 290 8167 416 8320
rect 482 8167 608 8320
rect 674 8167 800 8320
rect 866 8167 992 8320
rect 1058 8167 1184 8320
rect 1250 8167 1376 8320
rect 1828 8167 1860 8320
rect 1926 8167 2052 8320
rect 2118 8167 2244 8320
rect 2310 8167 2436 8320
rect 2502 8167 2628 8320
rect 2694 8167 2820 8320
rect 2886 8167 3012 8320
rect 3078 8167 3204 8320
rect 3656 8167 3688 8320
rect 3754 8167 3880 8320
rect 3946 8167 4072 8320
rect 4138 8167 4264 8320
rect 4330 8167 4456 8320
rect 4522 8167 4648 8320
rect 4714 8167 4840 8320
rect 4906 8167 5032 8320
rect 5484 8167 5516 8320
rect 5582 8167 5708 8320
rect 5774 8167 5900 8320
rect 5966 8167 6092 8320
rect 6158 8167 6284 8320
rect 6350 8167 6476 8320
rect 6542 8167 6668 8320
rect 6734 8167 6860 8320
rect 7312 8167 7344 8320
rect 7410 8167 7536 8320
rect 7602 8167 7728 8320
rect 7794 8167 7920 8320
rect 7986 8167 8112 8320
rect 8178 8167 8304 8320
rect 8370 8167 8496 8320
rect 8562 8167 8688 8320
rect 9140 8167 9172 8320
rect 9238 8167 9364 8320
rect 9430 8167 9556 8320
rect 9622 8167 9748 8320
rect 9814 8167 9940 8320
rect 10006 8167 10132 8320
rect 10198 8167 10324 8320
rect 10390 8167 10516 8320
rect 10968 8167 11000 8320
rect 11066 8167 11192 8320
rect 11258 8167 11384 8320
rect 11450 8167 11576 8320
rect 11642 8167 11768 8320
rect 11834 8167 11960 8320
rect 12026 8167 12152 8320
rect 12218 8167 12344 8320
rect 12796 8167 12828 8320
rect 12894 8167 13020 8320
rect 13086 8167 13212 8320
rect 13278 8167 13404 8320
rect 13470 8167 13596 8320
rect 13662 8167 13788 8320
rect 13854 8167 13980 8320
rect 14046 8167 14172 8320
rect 14624 8167 14656 8320
rect 14722 8167 14848 8320
rect 14914 8167 15040 8320
rect 15106 8167 15232 8320
rect 15298 8167 15424 8320
rect 15490 8167 15616 8320
rect 15682 8167 15808 8320
rect 15874 8167 16000 8320
rect 16452 8167 16484 8320
rect 16550 8167 16676 8320
rect 16742 8167 16868 8320
rect 16934 8167 17060 8320
rect 17126 8167 17252 8320
rect 17318 8167 17444 8320
rect 17510 8167 17636 8320
rect 17702 8167 17828 8320
rect 18280 8167 18312 8320
rect 18378 8167 18504 8320
rect 18570 8167 18696 8320
rect 18762 8167 18888 8320
rect 18954 8167 19080 8320
rect 19146 8167 19272 8320
rect 19338 8167 19464 8320
rect 19530 8167 19656 8320
rect 20108 8167 20140 8320
rect 20206 8167 20332 8320
rect 20398 8167 20524 8320
rect 20590 8167 20716 8320
rect 20782 8167 20908 8320
rect 20974 8167 21100 8320
rect 21166 8167 21292 8320
rect 21358 8167 21484 8320
rect 32 8157 98 8167
rect 224 8157 290 8167
rect 416 8157 482 8167
rect 608 8157 674 8167
rect 800 8157 866 8167
rect 992 8157 1058 8167
rect 1184 8157 1250 8167
rect 1376 8157 1442 8167
rect 1860 8157 1926 8167
rect 2052 8157 2118 8167
rect 2244 8157 2310 8167
rect 2436 8157 2502 8167
rect 2628 8157 2694 8167
rect 2820 8157 2886 8167
rect 3012 8157 3078 8167
rect 3204 8157 3270 8167
rect 3688 8157 3754 8167
rect 3880 8157 3946 8167
rect 4072 8157 4138 8167
rect 4264 8157 4330 8167
rect 4456 8157 4522 8167
rect 4648 8157 4714 8167
rect 4840 8157 4906 8167
rect 5032 8157 5098 8167
rect 5516 8157 5582 8167
rect 5708 8157 5774 8167
rect 5900 8157 5966 8167
rect 6092 8157 6158 8167
rect 6284 8157 6350 8167
rect 6476 8157 6542 8167
rect 6668 8157 6734 8167
rect 6860 8157 6926 8167
rect 7344 8157 7410 8167
rect 7536 8157 7602 8167
rect 7728 8157 7794 8167
rect 7920 8157 7986 8167
rect 8112 8157 8178 8167
rect 8304 8157 8370 8167
rect 8496 8157 8562 8167
rect 8688 8157 8754 8167
rect 9172 8157 9238 8167
rect 9364 8157 9430 8167
rect 9556 8157 9622 8167
rect 9748 8157 9814 8167
rect 9940 8157 10006 8167
rect 10132 8157 10198 8167
rect 10324 8157 10390 8167
rect 10516 8157 10582 8167
rect 11000 8157 11066 8167
rect 11192 8157 11258 8167
rect 11384 8157 11450 8167
rect 11576 8157 11642 8167
rect 11768 8157 11834 8167
rect 11960 8157 12026 8167
rect 12152 8157 12218 8167
rect 12344 8157 12410 8167
rect 12828 8157 12894 8167
rect 13020 8157 13086 8167
rect 13212 8157 13278 8167
rect 13404 8157 13470 8167
rect 13596 8157 13662 8167
rect 13788 8157 13854 8167
rect 13980 8157 14046 8167
rect 14172 8157 14238 8167
rect 14656 8157 14722 8167
rect 14848 8157 14914 8167
rect 15040 8157 15106 8167
rect 15232 8157 15298 8167
rect 15424 8157 15490 8167
rect 15616 8157 15682 8167
rect 15808 8157 15874 8167
rect 16000 8157 16066 8167
rect 16484 8157 16550 8167
rect 16676 8157 16742 8167
rect 16868 8157 16934 8167
rect 17060 8157 17126 8167
rect 17252 8157 17318 8167
rect 17444 8157 17510 8167
rect 17636 8157 17702 8167
rect 17828 8157 17894 8167
rect 18312 8157 18378 8167
rect 18504 8157 18570 8167
rect 18696 8157 18762 8167
rect 18888 8157 18954 8167
rect 19080 8157 19146 8167
rect 19272 8157 19338 8167
rect 19464 8157 19530 8167
rect 19656 8157 19722 8167
rect 20140 8157 20206 8167
rect 20332 8157 20398 8167
rect 20524 8157 20590 8167
rect 20716 8157 20782 8167
rect 20908 8157 20974 8167
rect 21100 8157 21166 8167
rect 21292 8157 21358 8167
rect 21484 8157 21550 8167
rect 128 8107 194 8117
rect 320 8107 386 8117
rect 512 8107 578 8117
rect 704 8107 770 8117
rect 896 8107 962 8117
rect 1088 8107 1154 8117
rect 1280 8107 1346 8117
rect 1472 8107 1528 8117
rect 1956 8107 2022 8117
rect 2148 8107 2214 8117
rect 2340 8107 2406 8117
rect 2532 8107 2598 8117
rect 2724 8107 2790 8117
rect 2916 8107 2982 8117
rect 3108 8107 3174 8117
rect 3300 8107 3356 8117
rect 3784 8107 3850 8117
rect 3976 8107 4042 8117
rect 4168 8107 4234 8117
rect 4360 8107 4426 8117
rect 4552 8107 4618 8117
rect 4744 8107 4810 8117
rect 4936 8107 5002 8117
rect 5128 8107 5184 8117
rect 5612 8107 5678 8117
rect 5804 8107 5870 8117
rect 5996 8107 6062 8117
rect 6188 8107 6254 8117
rect 6380 8107 6446 8117
rect 6572 8107 6638 8117
rect 6764 8107 6830 8117
rect 6956 8107 7012 8117
rect 7440 8107 7506 8117
rect 7632 8107 7698 8117
rect 7824 8107 7890 8117
rect 8016 8107 8082 8117
rect 8208 8107 8274 8117
rect 8400 8107 8466 8117
rect 8592 8107 8658 8117
rect 8784 8107 8840 8117
rect 9268 8107 9334 8117
rect 9460 8107 9526 8117
rect 9652 8107 9718 8117
rect 9844 8107 9910 8117
rect 10036 8107 10102 8117
rect 10228 8107 10294 8117
rect 10420 8107 10486 8117
rect 10612 8107 10668 8117
rect 11096 8107 11162 8117
rect 11288 8107 11354 8117
rect 11480 8107 11546 8117
rect 11672 8107 11738 8117
rect 11864 8107 11930 8117
rect 12056 8107 12122 8117
rect 12248 8107 12314 8117
rect 12440 8107 12496 8117
rect 12924 8107 12990 8117
rect 13116 8107 13182 8117
rect 13308 8107 13374 8117
rect 13500 8107 13566 8117
rect 13692 8107 13758 8117
rect 13884 8107 13950 8117
rect 14076 8107 14142 8117
rect 14268 8107 14324 8117
rect 14752 8107 14818 8117
rect 14944 8107 15010 8117
rect 15136 8107 15202 8117
rect 15328 8107 15394 8117
rect 15520 8107 15586 8117
rect 15712 8107 15778 8117
rect 15904 8107 15970 8117
rect 16096 8107 16152 8117
rect 16580 8107 16646 8117
rect 16772 8107 16838 8117
rect 16964 8107 17030 8117
rect 17156 8107 17222 8117
rect 17348 8107 17414 8117
rect 17540 8107 17606 8117
rect 17732 8107 17798 8117
rect 17924 8107 17980 8117
rect 18408 8107 18474 8117
rect 18600 8107 18666 8117
rect 18792 8107 18858 8117
rect 18984 8107 19050 8117
rect 19176 8107 19242 8117
rect 19368 8107 19434 8117
rect 19560 8107 19626 8117
rect 19752 8107 19808 8117
rect 20236 8107 20302 8117
rect 20428 8107 20494 8117
rect 20620 8107 20686 8117
rect 20812 8107 20878 8117
rect 21004 8107 21070 8117
rect 21196 8107 21262 8117
rect 21388 8107 21454 8117
rect 21580 8107 21636 8117
rect 0 7954 128 8107
rect 194 7954 320 8107
rect 386 7954 512 8107
rect 578 7954 704 8107
rect 770 7954 896 8107
rect 962 7954 1088 8107
rect 1154 7954 1280 8107
rect 1346 7954 1472 8107
rect 1528 7954 1708 8107
rect 1828 7954 1956 8107
rect 2022 7954 2148 8107
rect 2214 7954 2340 8107
rect 2406 7954 2532 8107
rect 2598 7954 2724 8107
rect 2790 7954 2916 8107
rect 2982 7954 3108 8107
rect 3174 7954 3300 8107
rect 3356 7954 3536 8107
rect 3656 7954 3784 8107
rect 3850 7954 3976 8107
rect 4042 7954 4168 8107
rect 4234 7954 4360 8107
rect 4426 7954 4552 8107
rect 4618 7954 4744 8107
rect 4810 7954 4936 8107
rect 5002 7954 5128 8107
rect 5184 7954 5364 8107
rect 5484 7954 5612 8107
rect 5678 7954 5804 8107
rect 5870 7954 5996 8107
rect 6062 7954 6188 8107
rect 6254 7954 6380 8107
rect 6446 7954 6572 8107
rect 6638 7954 6764 8107
rect 6830 7954 6956 8107
rect 7012 7954 7192 8107
rect 7312 7954 7440 8107
rect 7506 7954 7632 8107
rect 7698 7954 7824 8107
rect 7890 7954 8016 8107
rect 8082 7954 8208 8107
rect 8274 7954 8400 8107
rect 8466 7954 8592 8107
rect 8658 7954 8784 8107
rect 8840 7954 9020 8107
rect 9140 7954 9268 8107
rect 9334 7954 9460 8107
rect 9526 7954 9652 8107
rect 9718 7954 9844 8107
rect 9910 7954 10036 8107
rect 10102 7954 10228 8107
rect 10294 7954 10420 8107
rect 10486 7954 10612 8107
rect 10668 7954 10848 8107
rect 10968 7954 11096 8107
rect 11162 7954 11288 8107
rect 11354 7954 11480 8107
rect 11546 7954 11672 8107
rect 11738 7954 11864 8107
rect 11930 7954 12056 8107
rect 12122 7954 12248 8107
rect 12314 7954 12440 8107
rect 12496 7954 12676 8107
rect 12796 7954 12924 8107
rect 12990 7954 13116 8107
rect 13182 7954 13308 8107
rect 13374 7954 13500 8107
rect 13566 7954 13692 8107
rect 13758 7954 13884 8107
rect 13950 7954 14076 8107
rect 14142 7954 14268 8107
rect 14324 7954 14504 8107
rect 14624 7954 14752 8107
rect 14818 7954 14944 8107
rect 15010 7954 15136 8107
rect 15202 7954 15328 8107
rect 15394 7954 15520 8107
rect 15586 7954 15712 8107
rect 15778 7954 15904 8107
rect 15970 7954 16096 8107
rect 16152 7954 16332 8107
rect 16452 7954 16580 8107
rect 16646 7954 16772 8107
rect 16838 7954 16964 8107
rect 17030 7954 17156 8107
rect 17222 7954 17348 8107
rect 17414 7954 17540 8107
rect 17606 7954 17732 8107
rect 17798 7954 17924 8107
rect 17980 7954 18160 8107
rect 18280 7954 18408 8107
rect 18474 7954 18600 8107
rect 18666 7954 18792 8107
rect 18858 7954 18984 8107
rect 19050 7954 19176 8107
rect 19242 7954 19368 8107
rect 19434 7954 19560 8107
rect 19626 7954 19752 8107
rect 19808 7954 19988 8107
rect 20108 7954 20236 8107
rect 20302 7954 20428 8107
rect 20494 7954 20620 8107
rect 20686 7954 20812 8107
rect 20878 7954 21004 8107
rect 21070 7954 21196 8107
rect 21262 7954 21388 8107
rect 21454 7954 21580 8107
rect 21636 7954 21816 8107
rect 128 7944 194 7954
rect 320 7944 386 7954
rect 512 7944 578 7954
rect 704 7944 770 7954
rect 896 7944 962 7954
rect 1088 7944 1154 7954
rect 1280 7944 1346 7954
rect 1472 7944 1528 7954
rect 1956 7944 2022 7954
rect 2148 7944 2214 7954
rect 2340 7944 2406 7954
rect 2532 7944 2598 7954
rect 2724 7944 2790 7954
rect 2916 7944 2982 7954
rect 3108 7944 3174 7954
rect 3300 7944 3356 7954
rect 3784 7944 3850 7954
rect 3976 7944 4042 7954
rect 4168 7944 4234 7954
rect 4360 7944 4426 7954
rect 4552 7944 4618 7954
rect 4744 7944 4810 7954
rect 4936 7944 5002 7954
rect 5128 7944 5184 7954
rect 5612 7944 5678 7954
rect 5804 7944 5870 7954
rect 5996 7944 6062 7954
rect 6188 7944 6254 7954
rect 6380 7944 6446 7954
rect 6572 7944 6638 7954
rect 6764 7944 6830 7954
rect 6956 7944 7012 7954
rect 7440 7944 7506 7954
rect 7632 7944 7698 7954
rect 7824 7944 7890 7954
rect 8016 7944 8082 7954
rect 8208 7944 8274 7954
rect 8400 7944 8466 7954
rect 8592 7944 8658 7954
rect 8784 7944 8840 7954
rect 9268 7944 9334 7954
rect 9460 7944 9526 7954
rect 9652 7944 9718 7954
rect 9844 7944 9910 7954
rect 10036 7944 10102 7954
rect 10228 7944 10294 7954
rect 10420 7944 10486 7954
rect 10612 7944 10668 7954
rect 11096 7944 11162 7954
rect 11288 7944 11354 7954
rect 11480 7944 11546 7954
rect 11672 7944 11738 7954
rect 11864 7944 11930 7954
rect 12056 7944 12122 7954
rect 12248 7944 12314 7954
rect 12440 7944 12496 7954
rect 12924 7944 12990 7954
rect 13116 7944 13182 7954
rect 13308 7944 13374 7954
rect 13500 7944 13566 7954
rect 13692 7944 13758 7954
rect 13884 7944 13950 7954
rect 14076 7944 14142 7954
rect 14268 7944 14324 7954
rect 14752 7944 14818 7954
rect 14944 7944 15010 7954
rect 15136 7944 15202 7954
rect 15328 7944 15394 7954
rect 15520 7944 15586 7954
rect 15712 7944 15778 7954
rect 15904 7944 15970 7954
rect 16096 7944 16152 7954
rect 16580 7944 16646 7954
rect 16772 7944 16838 7954
rect 16964 7944 17030 7954
rect 17156 7944 17222 7954
rect 17348 7944 17414 7954
rect 17540 7944 17606 7954
rect 17732 7944 17798 7954
rect 17924 7944 17980 7954
rect 18408 7944 18474 7954
rect 18600 7944 18666 7954
rect 18792 7944 18858 7954
rect 18984 7944 19050 7954
rect 19176 7944 19242 7954
rect 19368 7944 19434 7954
rect 19560 7944 19626 7954
rect 19752 7944 19808 7954
rect 20236 7944 20302 7954
rect 20428 7944 20494 7954
rect 20620 7944 20686 7954
rect 20812 7944 20878 7954
rect 21004 7944 21070 7954
rect 21196 7944 21262 7954
rect 21388 7944 21454 7954
rect 21580 7944 21636 7954
rect 32 7606 98 7616
rect 224 7606 290 7616
rect 416 7606 482 7616
rect 608 7606 674 7616
rect 800 7606 866 7616
rect 992 7606 1058 7616
rect 1184 7606 1250 7616
rect 1376 7606 1442 7616
rect 1860 7606 1926 7616
rect 2052 7606 2118 7616
rect 2244 7606 2310 7616
rect 2436 7606 2502 7616
rect 2628 7606 2694 7616
rect 2820 7606 2886 7616
rect 3012 7606 3078 7616
rect 3204 7606 3270 7616
rect 3688 7606 3754 7616
rect 3880 7606 3946 7616
rect 4072 7606 4138 7616
rect 4264 7606 4330 7616
rect 4456 7606 4522 7616
rect 4648 7606 4714 7616
rect 4840 7606 4906 7616
rect 5032 7606 5098 7616
rect 5516 7606 5582 7616
rect 5708 7606 5774 7616
rect 5900 7606 5966 7616
rect 6092 7606 6158 7616
rect 6284 7606 6350 7616
rect 6476 7606 6542 7616
rect 6668 7606 6734 7616
rect 6860 7606 6926 7616
rect 7344 7606 7410 7616
rect 7536 7606 7602 7616
rect 7728 7606 7794 7616
rect 7920 7606 7986 7616
rect 8112 7606 8178 7616
rect 8304 7606 8370 7616
rect 8496 7606 8562 7616
rect 8688 7606 8754 7616
rect 9172 7606 9238 7616
rect 9364 7606 9430 7616
rect 9556 7606 9622 7616
rect 9748 7606 9814 7616
rect 9940 7606 10006 7616
rect 10132 7606 10198 7616
rect 10324 7606 10390 7616
rect 10516 7606 10582 7616
rect 11000 7606 11066 7616
rect 11192 7606 11258 7616
rect 11384 7606 11450 7616
rect 11576 7606 11642 7616
rect 11768 7606 11834 7616
rect 11960 7606 12026 7616
rect 12152 7606 12218 7616
rect 12344 7606 12410 7616
rect 12828 7606 12894 7616
rect 13020 7606 13086 7616
rect 13212 7606 13278 7616
rect 13404 7606 13470 7616
rect 13596 7606 13662 7616
rect 13788 7606 13854 7616
rect 13980 7606 14046 7616
rect 14172 7606 14238 7616
rect 14656 7606 14722 7616
rect 14848 7606 14914 7616
rect 15040 7606 15106 7616
rect 15232 7606 15298 7616
rect 15424 7606 15490 7616
rect 15616 7606 15682 7616
rect 15808 7606 15874 7616
rect 16000 7606 16066 7616
rect 16484 7606 16550 7616
rect 16676 7606 16742 7616
rect 16868 7606 16934 7616
rect 17060 7606 17126 7616
rect 17252 7606 17318 7616
rect 17444 7606 17510 7616
rect 17636 7606 17702 7616
rect 17828 7606 17894 7616
rect 18312 7606 18378 7616
rect 18504 7606 18570 7616
rect 18696 7606 18762 7616
rect 18888 7606 18954 7616
rect 19080 7606 19146 7616
rect 19272 7606 19338 7616
rect 19464 7606 19530 7616
rect 19656 7606 19722 7616
rect 20140 7606 20206 7616
rect 20332 7606 20398 7616
rect 20524 7606 20590 7616
rect 20716 7606 20782 7616
rect 20908 7606 20974 7616
rect 21100 7606 21166 7616
rect 21292 7606 21358 7616
rect 21484 7606 21550 7616
rect 0 7453 32 7606
rect 98 7453 224 7606
rect 290 7453 416 7606
rect 482 7453 608 7606
rect 674 7453 800 7606
rect 866 7453 992 7606
rect 1058 7453 1184 7606
rect 1250 7453 1376 7606
rect 1828 7453 1860 7606
rect 1926 7453 2052 7606
rect 2118 7453 2244 7606
rect 2310 7453 2436 7606
rect 2502 7453 2628 7606
rect 2694 7453 2820 7606
rect 2886 7453 3012 7606
rect 3078 7453 3204 7606
rect 3656 7453 3688 7606
rect 3754 7453 3880 7606
rect 3946 7453 4072 7606
rect 4138 7453 4264 7606
rect 4330 7453 4456 7606
rect 4522 7453 4648 7606
rect 4714 7453 4840 7606
rect 4906 7453 5032 7606
rect 5484 7453 5516 7606
rect 5582 7453 5708 7606
rect 5774 7453 5900 7606
rect 5966 7453 6092 7606
rect 6158 7453 6284 7606
rect 6350 7453 6476 7606
rect 6542 7453 6668 7606
rect 6734 7453 6860 7606
rect 7312 7453 7344 7606
rect 7410 7453 7536 7606
rect 7602 7453 7728 7606
rect 7794 7453 7920 7606
rect 7986 7453 8112 7606
rect 8178 7453 8304 7606
rect 8370 7453 8496 7606
rect 8562 7453 8688 7606
rect 9140 7453 9172 7606
rect 9238 7453 9364 7606
rect 9430 7453 9556 7606
rect 9622 7453 9748 7606
rect 9814 7453 9940 7606
rect 10006 7453 10132 7606
rect 10198 7453 10324 7606
rect 10390 7453 10516 7606
rect 10968 7453 11000 7606
rect 11066 7453 11192 7606
rect 11258 7453 11384 7606
rect 11450 7453 11576 7606
rect 11642 7453 11768 7606
rect 11834 7453 11960 7606
rect 12026 7453 12152 7606
rect 12218 7453 12344 7606
rect 12796 7453 12828 7606
rect 12894 7453 13020 7606
rect 13086 7453 13212 7606
rect 13278 7453 13404 7606
rect 13470 7453 13596 7606
rect 13662 7453 13788 7606
rect 13854 7453 13980 7606
rect 14046 7453 14172 7606
rect 14624 7453 14656 7606
rect 14722 7453 14848 7606
rect 14914 7453 15040 7606
rect 15106 7453 15232 7606
rect 15298 7453 15424 7606
rect 15490 7453 15616 7606
rect 15682 7453 15808 7606
rect 15874 7453 16000 7606
rect 16452 7453 16484 7606
rect 16550 7453 16676 7606
rect 16742 7453 16868 7606
rect 16934 7453 17060 7606
rect 17126 7453 17252 7606
rect 17318 7453 17444 7606
rect 17510 7453 17636 7606
rect 17702 7453 17828 7606
rect 18280 7453 18312 7606
rect 18378 7453 18504 7606
rect 18570 7453 18696 7606
rect 18762 7453 18888 7606
rect 18954 7453 19080 7606
rect 19146 7453 19272 7606
rect 19338 7453 19464 7606
rect 19530 7453 19656 7606
rect 20108 7453 20140 7606
rect 20206 7453 20332 7606
rect 20398 7453 20524 7606
rect 20590 7453 20716 7606
rect 20782 7453 20908 7606
rect 20974 7453 21100 7606
rect 21166 7453 21292 7606
rect 21358 7453 21484 7606
rect 32 7443 98 7453
rect 224 7443 290 7453
rect 416 7443 482 7453
rect 608 7443 674 7453
rect 800 7443 866 7453
rect 992 7443 1058 7453
rect 1184 7443 1250 7453
rect 1376 7443 1442 7453
rect 1860 7443 1926 7453
rect 2052 7443 2118 7453
rect 2244 7443 2310 7453
rect 2436 7443 2502 7453
rect 2628 7443 2694 7453
rect 2820 7443 2886 7453
rect 3012 7443 3078 7453
rect 3204 7443 3270 7453
rect 3688 7443 3754 7453
rect 3880 7443 3946 7453
rect 4072 7443 4138 7453
rect 4264 7443 4330 7453
rect 4456 7443 4522 7453
rect 4648 7443 4714 7453
rect 4840 7443 4906 7453
rect 5032 7443 5098 7453
rect 5516 7443 5582 7453
rect 5708 7443 5774 7453
rect 5900 7443 5966 7453
rect 6092 7443 6158 7453
rect 6284 7443 6350 7453
rect 6476 7443 6542 7453
rect 6668 7443 6734 7453
rect 6860 7443 6926 7453
rect 7344 7443 7410 7453
rect 7536 7443 7602 7453
rect 7728 7443 7794 7453
rect 7920 7443 7986 7453
rect 8112 7443 8178 7453
rect 8304 7443 8370 7453
rect 8496 7443 8562 7453
rect 8688 7443 8754 7453
rect 9172 7443 9238 7453
rect 9364 7443 9430 7453
rect 9556 7443 9622 7453
rect 9748 7443 9814 7453
rect 9940 7443 10006 7453
rect 10132 7443 10198 7453
rect 10324 7443 10390 7453
rect 10516 7443 10582 7453
rect 11000 7443 11066 7453
rect 11192 7443 11258 7453
rect 11384 7443 11450 7453
rect 11576 7443 11642 7453
rect 11768 7443 11834 7453
rect 11960 7443 12026 7453
rect 12152 7443 12218 7453
rect 12344 7443 12410 7453
rect 12828 7443 12894 7453
rect 13020 7443 13086 7453
rect 13212 7443 13278 7453
rect 13404 7443 13470 7453
rect 13596 7443 13662 7453
rect 13788 7443 13854 7453
rect 13980 7443 14046 7453
rect 14172 7443 14238 7453
rect 14656 7443 14722 7453
rect 14848 7443 14914 7453
rect 15040 7443 15106 7453
rect 15232 7443 15298 7453
rect 15424 7443 15490 7453
rect 15616 7443 15682 7453
rect 15808 7443 15874 7453
rect 16000 7443 16066 7453
rect 16484 7443 16550 7453
rect 16676 7443 16742 7453
rect 16868 7443 16934 7453
rect 17060 7443 17126 7453
rect 17252 7443 17318 7453
rect 17444 7443 17510 7453
rect 17636 7443 17702 7453
rect 17828 7443 17894 7453
rect 18312 7443 18378 7453
rect 18504 7443 18570 7453
rect 18696 7443 18762 7453
rect 18888 7443 18954 7453
rect 19080 7443 19146 7453
rect 19272 7443 19338 7453
rect 19464 7443 19530 7453
rect 19656 7443 19722 7453
rect 20140 7443 20206 7453
rect 20332 7443 20398 7453
rect 20524 7443 20590 7453
rect 20716 7443 20782 7453
rect 20908 7443 20974 7453
rect 21100 7443 21166 7453
rect 21292 7443 21358 7453
rect 21484 7443 21550 7453
rect 128 7393 194 7403
rect 320 7393 386 7403
rect 512 7393 578 7403
rect 704 7393 770 7403
rect 896 7393 962 7403
rect 1088 7393 1154 7403
rect 1280 7393 1346 7403
rect 1472 7393 1528 7403
rect 1956 7393 2022 7403
rect 2148 7393 2214 7403
rect 2340 7393 2406 7403
rect 2532 7393 2598 7403
rect 2724 7393 2790 7403
rect 2916 7393 2982 7403
rect 3108 7393 3174 7403
rect 3300 7393 3356 7403
rect 3784 7393 3850 7403
rect 3976 7393 4042 7403
rect 4168 7393 4234 7403
rect 4360 7393 4426 7403
rect 4552 7393 4618 7403
rect 4744 7393 4810 7403
rect 4936 7393 5002 7403
rect 5128 7393 5184 7403
rect 5612 7393 5678 7403
rect 5804 7393 5870 7403
rect 5996 7393 6062 7403
rect 6188 7393 6254 7403
rect 6380 7393 6446 7403
rect 6572 7393 6638 7403
rect 6764 7393 6830 7403
rect 6956 7393 7012 7403
rect 7440 7393 7506 7403
rect 7632 7393 7698 7403
rect 7824 7393 7890 7403
rect 8016 7393 8082 7403
rect 8208 7393 8274 7403
rect 8400 7393 8466 7403
rect 8592 7393 8658 7403
rect 8784 7393 8840 7403
rect 9268 7393 9334 7403
rect 9460 7393 9526 7403
rect 9652 7393 9718 7403
rect 9844 7393 9910 7403
rect 10036 7393 10102 7403
rect 10228 7393 10294 7403
rect 10420 7393 10486 7403
rect 10612 7393 10668 7403
rect 11096 7393 11162 7403
rect 11288 7393 11354 7403
rect 11480 7393 11546 7403
rect 11672 7393 11738 7403
rect 11864 7393 11930 7403
rect 12056 7393 12122 7403
rect 12248 7393 12314 7403
rect 12440 7393 12496 7403
rect 12924 7393 12990 7403
rect 13116 7393 13182 7403
rect 13308 7393 13374 7403
rect 13500 7393 13566 7403
rect 13692 7393 13758 7403
rect 13884 7393 13950 7403
rect 14076 7393 14142 7403
rect 14268 7393 14324 7403
rect 14752 7393 14818 7403
rect 14944 7393 15010 7403
rect 15136 7393 15202 7403
rect 15328 7393 15394 7403
rect 15520 7393 15586 7403
rect 15712 7393 15778 7403
rect 15904 7393 15970 7403
rect 16096 7393 16152 7403
rect 16580 7393 16646 7403
rect 16772 7393 16838 7403
rect 16964 7393 17030 7403
rect 17156 7393 17222 7403
rect 17348 7393 17414 7403
rect 17540 7393 17606 7403
rect 17732 7393 17798 7403
rect 17924 7393 17980 7403
rect 18408 7393 18474 7403
rect 18600 7393 18666 7403
rect 18792 7393 18858 7403
rect 18984 7393 19050 7403
rect 19176 7393 19242 7403
rect 19368 7393 19434 7403
rect 19560 7393 19626 7403
rect 19752 7393 19808 7403
rect 20236 7393 20302 7403
rect 20428 7393 20494 7403
rect 20620 7393 20686 7403
rect 20812 7393 20878 7403
rect 21004 7393 21070 7403
rect 21196 7393 21262 7403
rect 21388 7393 21454 7403
rect 21580 7393 21636 7403
rect 0 7240 128 7393
rect 194 7240 320 7393
rect 386 7240 512 7393
rect 578 7240 704 7393
rect 770 7240 896 7393
rect 962 7240 1088 7393
rect 1154 7240 1280 7393
rect 1346 7240 1472 7393
rect 1528 7240 1708 7393
rect 1828 7240 1956 7393
rect 2022 7240 2148 7393
rect 2214 7240 2340 7393
rect 2406 7240 2532 7393
rect 2598 7240 2724 7393
rect 2790 7240 2916 7393
rect 2982 7240 3108 7393
rect 3174 7240 3300 7393
rect 3356 7240 3536 7393
rect 3656 7240 3784 7393
rect 3850 7240 3976 7393
rect 4042 7240 4168 7393
rect 4234 7240 4360 7393
rect 4426 7240 4552 7393
rect 4618 7240 4744 7393
rect 4810 7240 4936 7393
rect 5002 7240 5128 7393
rect 5184 7240 5364 7393
rect 5484 7240 5612 7393
rect 5678 7240 5804 7393
rect 5870 7240 5996 7393
rect 6062 7240 6188 7393
rect 6254 7240 6380 7393
rect 6446 7240 6572 7393
rect 6638 7240 6764 7393
rect 6830 7240 6956 7393
rect 7012 7240 7192 7393
rect 7312 7240 7440 7393
rect 7506 7240 7632 7393
rect 7698 7240 7824 7393
rect 7890 7240 8016 7393
rect 8082 7240 8208 7393
rect 8274 7240 8400 7393
rect 8466 7240 8592 7393
rect 8658 7240 8784 7393
rect 8840 7240 9020 7393
rect 9140 7240 9268 7393
rect 9334 7240 9460 7393
rect 9526 7240 9652 7393
rect 9718 7240 9844 7393
rect 9910 7240 10036 7393
rect 10102 7240 10228 7393
rect 10294 7240 10420 7393
rect 10486 7240 10612 7393
rect 10668 7240 10848 7393
rect 10968 7240 11096 7393
rect 11162 7240 11288 7393
rect 11354 7240 11480 7393
rect 11546 7240 11672 7393
rect 11738 7240 11864 7393
rect 11930 7240 12056 7393
rect 12122 7240 12248 7393
rect 12314 7240 12440 7393
rect 12496 7240 12676 7393
rect 12796 7240 12924 7393
rect 12990 7240 13116 7393
rect 13182 7240 13308 7393
rect 13374 7240 13500 7393
rect 13566 7240 13692 7393
rect 13758 7240 13884 7393
rect 13950 7240 14076 7393
rect 14142 7240 14268 7393
rect 14324 7240 14504 7393
rect 14624 7240 14752 7393
rect 14818 7240 14944 7393
rect 15010 7240 15136 7393
rect 15202 7240 15328 7393
rect 15394 7240 15520 7393
rect 15586 7240 15712 7393
rect 15778 7240 15904 7393
rect 15970 7240 16096 7393
rect 16152 7240 16332 7393
rect 16452 7240 16580 7393
rect 16646 7240 16772 7393
rect 16838 7240 16964 7393
rect 17030 7240 17156 7393
rect 17222 7240 17348 7393
rect 17414 7240 17540 7393
rect 17606 7240 17732 7393
rect 17798 7240 17924 7393
rect 17980 7240 18160 7393
rect 18280 7240 18408 7393
rect 18474 7240 18600 7393
rect 18666 7240 18792 7393
rect 18858 7240 18984 7393
rect 19050 7240 19176 7393
rect 19242 7240 19368 7393
rect 19434 7240 19560 7393
rect 19626 7240 19752 7393
rect 19808 7240 19988 7393
rect 20108 7240 20236 7393
rect 20302 7240 20428 7393
rect 20494 7240 20620 7393
rect 20686 7240 20812 7393
rect 20878 7240 21004 7393
rect 21070 7240 21196 7393
rect 21262 7240 21388 7393
rect 21454 7240 21580 7393
rect 21636 7240 21816 7393
rect 128 7230 194 7240
rect 320 7230 386 7240
rect 512 7230 578 7240
rect 704 7230 770 7240
rect 896 7230 962 7240
rect 1088 7230 1154 7240
rect 1280 7230 1346 7240
rect 1472 7230 1528 7240
rect 1956 7230 2022 7240
rect 2148 7230 2214 7240
rect 2340 7230 2406 7240
rect 2532 7230 2598 7240
rect 2724 7230 2790 7240
rect 2916 7230 2982 7240
rect 3108 7230 3174 7240
rect 3300 7230 3356 7240
rect 3784 7230 3850 7240
rect 3976 7230 4042 7240
rect 4168 7230 4234 7240
rect 4360 7230 4426 7240
rect 4552 7230 4618 7240
rect 4744 7230 4810 7240
rect 4936 7230 5002 7240
rect 5128 7230 5184 7240
rect 5612 7230 5678 7240
rect 5804 7230 5870 7240
rect 5996 7230 6062 7240
rect 6188 7230 6254 7240
rect 6380 7230 6446 7240
rect 6572 7230 6638 7240
rect 6764 7230 6830 7240
rect 6956 7230 7012 7240
rect 7440 7230 7506 7240
rect 7632 7230 7698 7240
rect 7824 7230 7890 7240
rect 8016 7230 8082 7240
rect 8208 7230 8274 7240
rect 8400 7230 8466 7240
rect 8592 7230 8658 7240
rect 8784 7230 8840 7240
rect 9268 7230 9334 7240
rect 9460 7230 9526 7240
rect 9652 7230 9718 7240
rect 9844 7230 9910 7240
rect 10036 7230 10102 7240
rect 10228 7230 10294 7240
rect 10420 7230 10486 7240
rect 10612 7230 10668 7240
rect 11096 7230 11162 7240
rect 11288 7230 11354 7240
rect 11480 7230 11546 7240
rect 11672 7230 11738 7240
rect 11864 7230 11930 7240
rect 12056 7230 12122 7240
rect 12248 7230 12314 7240
rect 12440 7230 12496 7240
rect 12924 7230 12990 7240
rect 13116 7230 13182 7240
rect 13308 7230 13374 7240
rect 13500 7230 13566 7240
rect 13692 7230 13758 7240
rect 13884 7230 13950 7240
rect 14076 7230 14142 7240
rect 14268 7230 14324 7240
rect 14752 7230 14818 7240
rect 14944 7230 15010 7240
rect 15136 7230 15202 7240
rect 15328 7230 15394 7240
rect 15520 7230 15586 7240
rect 15712 7230 15778 7240
rect 15904 7230 15970 7240
rect 16096 7230 16152 7240
rect 16580 7230 16646 7240
rect 16772 7230 16838 7240
rect 16964 7230 17030 7240
rect 17156 7230 17222 7240
rect 17348 7230 17414 7240
rect 17540 7230 17606 7240
rect 17732 7230 17798 7240
rect 17924 7230 17980 7240
rect 18408 7230 18474 7240
rect 18600 7230 18666 7240
rect 18792 7230 18858 7240
rect 18984 7230 19050 7240
rect 19176 7230 19242 7240
rect 19368 7230 19434 7240
rect 19560 7230 19626 7240
rect 19752 7230 19808 7240
rect 20236 7230 20302 7240
rect 20428 7230 20494 7240
rect 20620 7230 20686 7240
rect 20812 7230 20878 7240
rect 21004 7230 21070 7240
rect 21196 7230 21262 7240
rect 21388 7230 21454 7240
rect 21580 7230 21636 7240
rect 32 6892 98 6902
rect 224 6892 290 6902
rect 416 6892 482 6902
rect 608 6892 674 6902
rect 800 6892 866 6902
rect 992 6892 1058 6902
rect 1184 6892 1250 6902
rect 1376 6892 1442 6902
rect 1860 6892 1926 6902
rect 2052 6892 2118 6902
rect 2244 6892 2310 6902
rect 2436 6892 2502 6902
rect 2628 6892 2694 6902
rect 2820 6892 2886 6902
rect 3012 6892 3078 6902
rect 3204 6892 3270 6902
rect 3688 6892 3754 6902
rect 3880 6892 3946 6902
rect 4072 6892 4138 6902
rect 4264 6892 4330 6902
rect 4456 6892 4522 6902
rect 4648 6892 4714 6902
rect 4840 6892 4906 6902
rect 5032 6892 5098 6902
rect 5516 6892 5582 6902
rect 5708 6892 5774 6902
rect 5900 6892 5966 6902
rect 6092 6892 6158 6902
rect 6284 6892 6350 6902
rect 6476 6892 6542 6902
rect 6668 6892 6734 6902
rect 6860 6892 6926 6902
rect 7344 6892 7410 6902
rect 7536 6892 7602 6902
rect 7728 6892 7794 6902
rect 7920 6892 7986 6902
rect 8112 6892 8178 6902
rect 8304 6892 8370 6902
rect 8496 6892 8562 6902
rect 8688 6892 8754 6902
rect 9172 6892 9238 6902
rect 9364 6892 9430 6902
rect 9556 6892 9622 6902
rect 9748 6892 9814 6902
rect 9940 6892 10006 6902
rect 10132 6892 10198 6902
rect 10324 6892 10390 6902
rect 10516 6892 10582 6902
rect 11000 6892 11066 6902
rect 11192 6892 11258 6902
rect 11384 6892 11450 6902
rect 11576 6892 11642 6902
rect 11768 6892 11834 6902
rect 11960 6892 12026 6902
rect 12152 6892 12218 6902
rect 12344 6892 12410 6902
rect 12828 6892 12894 6902
rect 13020 6892 13086 6902
rect 13212 6892 13278 6902
rect 13404 6892 13470 6902
rect 13596 6892 13662 6902
rect 13788 6892 13854 6902
rect 13980 6892 14046 6902
rect 14172 6892 14238 6902
rect 14656 6892 14722 6902
rect 14848 6892 14914 6902
rect 15040 6892 15106 6902
rect 15232 6892 15298 6902
rect 15424 6892 15490 6902
rect 15616 6892 15682 6902
rect 15808 6892 15874 6902
rect 16000 6892 16066 6902
rect 16484 6892 16550 6902
rect 16676 6892 16742 6902
rect 16868 6892 16934 6902
rect 17060 6892 17126 6902
rect 17252 6892 17318 6902
rect 17444 6892 17510 6902
rect 17636 6892 17702 6902
rect 17828 6892 17894 6902
rect 18312 6892 18378 6902
rect 18504 6892 18570 6902
rect 18696 6892 18762 6902
rect 18888 6892 18954 6902
rect 19080 6892 19146 6902
rect 19272 6892 19338 6902
rect 19464 6892 19530 6902
rect 19656 6892 19722 6902
rect 20140 6892 20206 6902
rect 20332 6892 20398 6902
rect 20524 6892 20590 6902
rect 20716 6892 20782 6902
rect 20908 6892 20974 6902
rect 21100 6892 21166 6902
rect 21292 6892 21358 6902
rect 21484 6892 21550 6902
rect 0 6739 32 6892
rect 98 6739 224 6892
rect 290 6739 416 6892
rect 482 6739 608 6892
rect 674 6739 800 6892
rect 866 6739 992 6892
rect 1058 6739 1184 6892
rect 1250 6739 1376 6892
rect 1828 6739 1860 6892
rect 1926 6739 2052 6892
rect 2118 6739 2244 6892
rect 2310 6739 2436 6892
rect 2502 6739 2628 6892
rect 2694 6739 2820 6892
rect 2886 6739 3012 6892
rect 3078 6739 3204 6892
rect 3656 6739 3688 6892
rect 3754 6739 3880 6892
rect 3946 6739 4072 6892
rect 4138 6739 4264 6892
rect 4330 6739 4456 6892
rect 4522 6739 4648 6892
rect 4714 6739 4840 6892
rect 4906 6739 5032 6892
rect 5484 6739 5516 6892
rect 5582 6739 5708 6892
rect 5774 6739 5900 6892
rect 5966 6739 6092 6892
rect 6158 6739 6284 6892
rect 6350 6739 6476 6892
rect 6542 6739 6668 6892
rect 6734 6739 6860 6892
rect 7312 6739 7344 6892
rect 7410 6739 7536 6892
rect 7602 6739 7728 6892
rect 7794 6739 7920 6892
rect 7986 6739 8112 6892
rect 8178 6739 8304 6892
rect 8370 6739 8496 6892
rect 8562 6739 8688 6892
rect 9140 6739 9172 6892
rect 9238 6739 9364 6892
rect 9430 6739 9556 6892
rect 9622 6739 9748 6892
rect 9814 6739 9940 6892
rect 10006 6739 10132 6892
rect 10198 6739 10324 6892
rect 10390 6739 10516 6892
rect 10968 6739 11000 6892
rect 11066 6739 11192 6892
rect 11258 6739 11384 6892
rect 11450 6739 11576 6892
rect 11642 6739 11768 6892
rect 11834 6739 11960 6892
rect 12026 6739 12152 6892
rect 12218 6739 12344 6892
rect 12796 6739 12828 6892
rect 12894 6739 13020 6892
rect 13086 6739 13212 6892
rect 13278 6739 13404 6892
rect 13470 6739 13596 6892
rect 13662 6739 13788 6892
rect 13854 6739 13980 6892
rect 14046 6739 14172 6892
rect 14624 6739 14656 6892
rect 14722 6739 14848 6892
rect 14914 6739 15040 6892
rect 15106 6739 15232 6892
rect 15298 6739 15424 6892
rect 15490 6739 15616 6892
rect 15682 6739 15808 6892
rect 15874 6739 16000 6892
rect 16452 6739 16484 6892
rect 16550 6739 16676 6892
rect 16742 6739 16868 6892
rect 16934 6739 17060 6892
rect 17126 6739 17252 6892
rect 17318 6739 17444 6892
rect 17510 6739 17636 6892
rect 17702 6739 17828 6892
rect 18280 6739 18312 6892
rect 18378 6739 18504 6892
rect 18570 6739 18696 6892
rect 18762 6739 18888 6892
rect 18954 6739 19080 6892
rect 19146 6739 19272 6892
rect 19338 6739 19464 6892
rect 19530 6739 19656 6892
rect 20108 6739 20140 6892
rect 20206 6739 20332 6892
rect 20398 6739 20524 6892
rect 20590 6739 20716 6892
rect 20782 6739 20908 6892
rect 20974 6739 21100 6892
rect 21166 6739 21292 6892
rect 21358 6739 21484 6892
rect 32 6729 98 6739
rect 224 6729 290 6739
rect 416 6729 482 6739
rect 608 6729 674 6739
rect 800 6729 866 6739
rect 992 6729 1058 6739
rect 1184 6729 1250 6739
rect 1376 6729 1442 6739
rect 1860 6729 1926 6739
rect 2052 6729 2118 6739
rect 2244 6729 2310 6739
rect 2436 6729 2502 6739
rect 2628 6729 2694 6739
rect 2820 6729 2886 6739
rect 3012 6729 3078 6739
rect 3204 6729 3270 6739
rect 3688 6729 3754 6739
rect 3880 6729 3946 6739
rect 4072 6729 4138 6739
rect 4264 6729 4330 6739
rect 4456 6729 4522 6739
rect 4648 6729 4714 6739
rect 4840 6729 4906 6739
rect 5032 6729 5098 6739
rect 5516 6729 5582 6739
rect 5708 6729 5774 6739
rect 5900 6729 5966 6739
rect 6092 6729 6158 6739
rect 6284 6729 6350 6739
rect 6476 6729 6542 6739
rect 6668 6729 6734 6739
rect 6860 6729 6926 6739
rect 7344 6729 7410 6739
rect 7536 6729 7602 6739
rect 7728 6729 7794 6739
rect 7920 6729 7986 6739
rect 8112 6729 8178 6739
rect 8304 6729 8370 6739
rect 8496 6729 8562 6739
rect 8688 6729 8754 6739
rect 9172 6729 9238 6739
rect 9364 6729 9430 6739
rect 9556 6729 9622 6739
rect 9748 6729 9814 6739
rect 9940 6729 10006 6739
rect 10132 6729 10198 6739
rect 10324 6729 10390 6739
rect 10516 6729 10582 6739
rect 11000 6729 11066 6739
rect 11192 6729 11258 6739
rect 11384 6729 11450 6739
rect 11576 6729 11642 6739
rect 11768 6729 11834 6739
rect 11960 6729 12026 6739
rect 12152 6729 12218 6739
rect 12344 6729 12410 6739
rect 12828 6729 12894 6739
rect 13020 6729 13086 6739
rect 13212 6729 13278 6739
rect 13404 6729 13470 6739
rect 13596 6729 13662 6739
rect 13788 6729 13854 6739
rect 13980 6729 14046 6739
rect 14172 6729 14238 6739
rect 14656 6729 14722 6739
rect 14848 6729 14914 6739
rect 15040 6729 15106 6739
rect 15232 6729 15298 6739
rect 15424 6729 15490 6739
rect 15616 6729 15682 6739
rect 15808 6729 15874 6739
rect 16000 6729 16066 6739
rect 16484 6729 16550 6739
rect 16676 6729 16742 6739
rect 16868 6729 16934 6739
rect 17060 6729 17126 6739
rect 17252 6729 17318 6739
rect 17444 6729 17510 6739
rect 17636 6729 17702 6739
rect 17828 6729 17894 6739
rect 18312 6729 18378 6739
rect 18504 6729 18570 6739
rect 18696 6729 18762 6739
rect 18888 6729 18954 6739
rect 19080 6729 19146 6739
rect 19272 6729 19338 6739
rect 19464 6729 19530 6739
rect 19656 6729 19722 6739
rect 20140 6729 20206 6739
rect 20332 6729 20398 6739
rect 20524 6729 20590 6739
rect 20716 6729 20782 6739
rect 20908 6729 20974 6739
rect 21100 6729 21166 6739
rect 21292 6729 21358 6739
rect 21484 6729 21550 6739
rect 128 6679 194 6689
rect 320 6679 386 6689
rect 512 6679 578 6689
rect 704 6679 770 6689
rect 896 6679 962 6689
rect 1088 6679 1154 6689
rect 1280 6679 1346 6689
rect 1472 6679 1528 6689
rect 1956 6679 2022 6689
rect 2148 6679 2214 6689
rect 2340 6679 2406 6689
rect 2532 6679 2598 6689
rect 2724 6679 2790 6689
rect 2916 6679 2982 6689
rect 3108 6679 3174 6689
rect 3300 6679 3356 6689
rect 3784 6679 3850 6689
rect 3976 6679 4042 6689
rect 4168 6679 4234 6689
rect 4360 6679 4426 6689
rect 4552 6679 4618 6689
rect 4744 6679 4810 6689
rect 4936 6679 5002 6689
rect 5128 6679 5184 6689
rect 5612 6679 5678 6689
rect 5804 6679 5870 6689
rect 5996 6679 6062 6689
rect 6188 6679 6254 6689
rect 6380 6679 6446 6689
rect 6572 6679 6638 6689
rect 6764 6679 6830 6689
rect 6956 6679 7012 6689
rect 7440 6679 7506 6689
rect 7632 6679 7698 6689
rect 7824 6679 7890 6689
rect 8016 6679 8082 6689
rect 8208 6679 8274 6689
rect 8400 6679 8466 6689
rect 8592 6679 8658 6689
rect 8784 6679 8840 6689
rect 9268 6679 9334 6689
rect 9460 6679 9526 6689
rect 9652 6679 9718 6689
rect 9844 6679 9910 6689
rect 10036 6679 10102 6689
rect 10228 6679 10294 6689
rect 10420 6679 10486 6689
rect 10612 6679 10668 6689
rect 11096 6679 11162 6689
rect 11288 6679 11354 6689
rect 11480 6679 11546 6689
rect 11672 6679 11738 6689
rect 11864 6679 11930 6689
rect 12056 6679 12122 6689
rect 12248 6679 12314 6689
rect 12440 6679 12496 6689
rect 12924 6679 12990 6689
rect 13116 6679 13182 6689
rect 13308 6679 13374 6689
rect 13500 6679 13566 6689
rect 13692 6679 13758 6689
rect 13884 6679 13950 6689
rect 14076 6679 14142 6689
rect 14268 6679 14324 6689
rect 14752 6679 14818 6689
rect 14944 6679 15010 6689
rect 15136 6679 15202 6689
rect 15328 6679 15394 6689
rect 15520 6679 15586 6689
rect 15712 6679 15778 6689
rect 15904 6679 15970 6689
rect 16096 6679 16152 6689
rect 16580 6679 16646 6689
rect 16772 6679 16838 6689
rect 16964 6679 17030 6689
rect 17156 6679 17222 6689
rect 17348 6679 17414 6689
rect 17540 6679 17606 6689
rect 17732 6679 17798 6689
rect 17924 6679 17980 6689
rect 18408 6679 18474 6689
rect 18600 6679 18666 6689
rect 18792 6679 18858 6689
rect 18984 6679 19050 6689
rect 19176 6679 19242 6689
rect 19368 6679 19434 6689
rect 19560 6679 19626 6689
rect 19752 6679 19808 6689
rect 20236 6679 20302 6689
rect 20428 6679 20494 6689
rect 20620 6679 20686 6689
rect 20812 6679 20878 6689
rect 21004 6679 21070 6689
rect 21196 6679 21262 6689
rect 21388 6679 21454 6689
rect 21580 6679 21636 6689
rect 0 6526 128 6679
rect 194 6526 320 6679
rect 386 6526 512 6679
rect 578 6526 704 6679
rect 770 6526 896 6679
rect 962 6526 1088 6679
rect 1154 6526 1280 6679
rect 1346 6526 1472 6679
rect 1528 6526 1708 6679
rect 1828 6526 1956 6679
rect 2022 6526 2148 6679
rect 2214 6526 2340 6679
rect 2406 6526 2532 6679
rect 2598 6526 2724 6679
rect 2790 6526 2916 6679
rect 2982 6526 3108 6679
rect 3174 6526 3300 6679
rect 3356 6526 3536 6679
rect 3656 6526 3784 6679
rect 3850 6526 3976 6679
rect 4042 6526 4168 6679
rect 4234 6526 4360 6679
rect 4426 6526 4552 6679
rect 4618 6526 4744 6679
rect 4810 6526 4936 6679
rect 5002 6526 5128 6679
rect 5184 6526 5364 6679
rect 5484 6526 5612 6679
rect 5678 6526 5804 6679
rect 5870 6526 5996 6679
rect 6062 6526 6188 6679
rect 6254 6526 6380 6679
rect 6446 6526 6572 6679
rect 6638 6526 6764 6679
rect 6830 6526 6956 6679
rect 7012 6526 7192 6679
rect 7312 6526 7440 6679
rect 7506 6526 7632 6679
rect 7698 6526 7824 6679
rect 7890 6526 8016 6679
rect 8082 6526 8208 6679
rect 8274 6526 8400 6679
rect 8466 6526 8592 6679
rect 8658 6526 8784 6679
rect 8840 6526 9020 6679
rect 9140 6526 9268 6679
rect 9334 6526 9460 6679
rect 9526 6526 9652 6679
rect 9718 6526 9844 6679
rect 9910 6526 10036 6679
rect 10102 6526 10228 6679
rect 10294 6526 10420 6679
rect 10486 6526 10612 6679
rect 10668 6526 10848 6679
rect 10968 6526 11096 6679
rect 11162 6526 11288 6679
rect 11354 6526 11480 6679
rect 11546 6526 11672 6679
rect 11738 6526 11864 6679
rect 11930 6526 12056 6679
rect 12122 6526 12248 6679
rect 12314 6526 12440 6679
rect 12496 6526 12676 6679
rect 12796 6526 12924 6679
rect 12990 6526 13116 6679
rect 13182 6526 13308 6679
rect 13374 6526 13500 6679
rect 13566 6526 13692 6679
rect 13758 6526 13884 6679
rect 13950 6526 14076 6679
rect 14142 6526 14268 6679
rect 14324 6526 14504 6679
rect 14624 6526 14752 6679
rect 14818 6526 14944 6679
rect 15010 6526 15136 6679
rect 15202 6526 15328 6679
rect 15394 6526 15520 6679
rect 15586 6526 15712 6679
rect 15778 6526 15904 6679
rect 15970 6526 16096 6679
rect 16152 6526 16332 6679
rect 16452 6526 16580 6679
rect 16646 6526 16772 6679
rect 16838 6526 16964 6679
rect 17030 6526 17156 6679
rect 17222 6526 17348 6679
rect 17414 6526 17540 6679
rect 17606 6526 17732 6679
rect 17798 6526 17924 6679
rect 17980 6526 18160 6679
rect 18280 6526 18408 6679
rect 18474 6526 18600 6679
rect 18666 6526 18792 6679
rect 18858 6526 18984 6679
rect 19050 6526 19176 6679
rect 19242 6526 19368 6679
rect 19434 6526 19560 6679
rect 19626 6526 19752 6679
rect 19808 6526 19988 6679
rect 20108 6526 20236 6679
rect 20302 6526 20428 6679
rect 20494 6526 20620 6679
rect 20686 6526 20812 6679
rect 20878 6526 21004 6679
rect 21070 6526 21196 6679
rect 21262 6526 21388 6679
rect 21454 6526 21580 6679
rect 21636 6526 21816 6679
rect 128 6516 194 6526
rect 320 6516 386 6526
rect 512 6516 578 6526
rect 704 6516 770 6526
rect 896 6516 962 6526
rect 1088 6516 1154 6526
rect 1280 6516 1346 6526
rect 1472 6516 1528 6526
rect 1956 6516 2022 6526
rect 2148 6516 2214 6526
rect 2340 6516 2406 6526
rect 2532 6516 2598 6526
rect 2724 6516 2790 6526
rect 2916 6516 2982 6526
rect 3108 6516 3174 6526
rect 3300 6516 3356 6526
rect 3784 6516 3850 6526
rect 3976 6516 4042 6526
rect 4168 6516 4234 6526
rect 4360 6516 4426 6526
rect 4552 6516 4618 6526
rect 4744 6516 4810 6526
rect 4936 6516 5002 6526
rect 5128 6516 5184 6526
rect 5612 6516 5678 6526
rect 5804 6516 5870 6526
rect 5996 6516 6062 6526
rect 6188 6516 6254 6526
rect 6380 6516 6446 6526
rect 6572 6516 6638 6526
rect 6764 6516 6830 6526
rect 6956 6516 7012 6526
rect 7440 6516 7506 6526
rect 7632 6516 7698 6526
rect 7824 6516 7890 6526
rect 8016 6516 8082 6526
rect 8208 6516 8274 6526
rect 8400 6516 8466 6526
rect 8592 6516 8658 6526
rect 8784 6516 8840 6526
rect 9268 6516 9334 6526
rect 9460 6516 9526 6526
rect 9652 6516 9718 6526
rect 9844 6516 9910 6526
rect 10036 6516 10102 6526
rect 10228 6516 10294 6526
rect 10420 6516 10486 6526
rect 10612 6516 10668 6526
rect 11096 6516 11162 6526
rect 11288 6516 11354 6526
rect 11480 6516 11546 6526
rect 11672 6516 11738 6526
rect 11864 6516 11930 6526
rect 12056 6516 12122 6526
rect 12248 6516 12314 6526
rect 12440 6516 12496 6526
rect 12924 6516 12990 6526
rect 13116 6516 13182 6526
rect 13308 6516 13374 6526
rect 13500 6516 13566 6526
rect 13692 6516 13758 6526
rect 13884 6516 13950 6526
rect 14076 6516 14142 6526
rect 14268 6516 14324 6526
rect 14752 6516 14818 6526
rect 14944 6516 15010 6526
rect 15136 6516 15202 6526
rect 15328 6516 15394 6526
rect 15520 6516 15586 6526
rect 15712 6516 15778 6526
rect 15904 6516 15970 6526
rect 16096 6516 16152 6526
rect 16580 6516 16646 6526
rect 16772 6516 16838 6526
rect 16964 6516 17030 6526
rect 17156 6516 17222 6526
rect 17348 6516 17414 6526
rect 17540 6516 17606 6526
rect 17732 6516 17798 6526
rect 17924 6516 17980 6526
rect 18408 6516 18474 6526
rect 18600 6516 18666 6526
rect 18792 6516 18858 6526
rect 18984 6516 19050 6526
rect 19176 6516 19242 6526
rect 19368 6516 19434 6526
rect 19560 6516 19626 6526
rect 19752 6516 19808 6526
rect 20236 6516 20302 6526
rect 20428 6516 20494 6526
rect 20620 6516 20686 6526
rect 20812 6516 20878 6526
rect 21004 6516 21070 6526
rect 21196 6516 21262 6526
rect 21388 6516 21454 6526
rect 21580 6516 21636 6526
rect 32 6178 98 6188
rect 224 6178 290 6188
rect 416 6178 482 6188
rect 608 6178 674 6188
rect 800 6178 866 6188
rect 992 6178 1058 6188
rect 1184 6178 1250 6188
rect 1376 6178 1442 6188
rect 1860 6178 1926 6188
rect 2052 6178 2118 6188
rect 2244 6178 2310 6188
rect 2436 6178 2502 6188
rect 2628 6178 2694 6188
rect 2820 6178 2886 6188
rect 3012 6178 3078 6188
rect 3204 6178 3270 6188
rect 3688 6178 3754 6188
rect 3880 6178 3946 6188
rect 4072 6178 4138 6188
rect 4264 6178 4330 6188
rect 4456 6178 4522 6188
rect 4648 6178 4714 6188
rect 4840 6178 4906 6188
rect 5032 6178 5098 6188
rect 5516 6178 5582 6188
rect 5708 6178 5774 6188
rect 5900 6178 5966 6188
rect 6092 6178 6158 6188
rect 6284 6178 6350 6188
rect 6476 6178 6542 6188
rect 6668 6178 6734 6188
rect 6860 6178 6926 6188
rect 7344 6178 7410 6188
rect 7536 6178 7602 6188
rect 7728 6178 7794 6188
rect 7920 6178 7986 6188
rect 8112 6178 8178 6188
rect 8304 6178 8370 6188
rect 8496 6178 8562 6188
rect 8688 6178 8754 6188
rect 9172 6178 9238 6188
rect 9364 6178 9430 6188
rect 9556 6178 9622 6188
rect 9748 6178 9814 6188
rect 9940 6178 10006 6188
rect 10132 6178 10198 6188
rect 10324 6178 10390 6188
rect 10516 6178 10582 6188
rect 11000 6178 11066 6188
rect 11192 6178 11258 6188
rect 11384 6178 11450 6188
rect 11576 6178 11642 6188
rect 11768 6178 11834 6188
rect 11960 6178 12026 6188
rect 12152 6178 12218 6188
rect 12344 6178 12410 6188
rect 12828 6178 12894 6188
rect 13020 6178 13086 6188
rect 13212 6178 13278 6188
rect 13404 6178 13470 6188
rect 13596 6178 13662 6188
rect 13788 6178 13854 6188
rect 13980 6178 14046 6188
rect 14172 6178 14238 6188
rect 14656 6178 14722 6188
rect 14848 6178 14914 6188
rect 15040 6178 15106 6188
rect 15232 6178 15298 6188
rect 15424 6178 15490 6188
rect 15616 6178 15682 6188
rect 15808 6178 15874 6188
rect 16000 6178 16066 6188
rect 16484 6178 16550 6188
rect 16676 6178 16742 6188
rect 16868 6178 16934 6188
rect 17060 6178 17126 6188
rect 17252 6178 17318 6188
rect 17444 6178 17510 6188
rect 17636 6178 17702 6188
rect 17828 6178 17894 6188
rect 18312 6178 18378 6188
rect 18504 6178 18570 6188
rect 18696 6178 18762 6188
rect 18888 6178 18954 6188
rect 19080 6178 19146 6188
rect 19272 6178 19338 6188
rect 19464 6178 19530 6188
rect 19656 6178 19722 6188
rect 20140 6178 20206 6188
rect 20332 6178 20398 6188
rect 20524 6178 20590 6188
rect 20716 6178 20782 6188
rect 20908 6178 20974 6188
rect 21100 6178 21166 6188
rect 21292 6178 21358 6188
rect 21484 6178 21550 6188
rect 0 6025 32 6178
rect 98 6025 224 6178
rect 290 6025 416 6178
rect 482 6025 608 6178
rect 674 6025 800 6178
rect 866 6025 992 6178
rect 1058 6025 1184 6178
rect 1250 6025 1376 6178
rect 1828 6025 1860 6178
rect 1926 6025 2052 6178
rect 2118 6025 2244 6178
rect 2310 6025 2436 6178
rect 2502 6025 2628 6178
rect 2694 6025 2820 6178
rect 2886 6025 3012 6178
rect 3078 6025 3204 6178
rect 3656 6025 3688 6178
rect 3754 6025 3880 6178
rect 3946 6025 4072 6178
rect 4138 6025 4264 6178
rect 4330 6025 4456 6178
rect 4522 6025 4648 6178
rect 4714 6025 4840 6178
rect 4906 6025 5032 6178
rect 5484 6025 5516 6178
rect 5582 6025 5708 6178
rect 5774 6025 5900 6178
rect 5966 6025 6092 6178
rect 6158 6025 6284 6178
rect 6350 6025 6476 6178
rect 6542 6025 6668 6178
rect 6734 6025 6860 6178
rect 7312 6025 7344 6178
rect 7410 6025 7536 6178
rect 7602 6025 7728 6178
rect 7794 6025 7920 6178
rect 7986 6025 8112 6178
rect 8178 6025 8304 6178
rect 8370 6025 8496 6178
rect 8562 6025 8688 6178
rect 9140 6025 9172 6178
rect 9238 6025 9364 6178
rect 9430 6025 9556 6178
rect 9622 6025 9748 6178
rect 9814 6025 9940 6178
rect 10006 6025 10132 6178
rect 10198 6025 10324 6178
rect 10390 6025 10516 6178
rect 10968 6025 11000 6178
rect 11066 6025 11192 6178
rect 11258 6025 11384 6178
rect 11450 6025 11576 6178
rect 11642 6025 11768 6178
rect 11834 6025 11960 6178
rect 12026 6025 12152 6178
rect 12218 6025 12344 6178
rect 12796 6025 12828 6178
rect 12894 6025 13020 6178
rect 13086 6025 13212 6178
rect 13278 6025 13404 6178
rect 13470 6025 13596 6178
rect 13662 6025 13788 6178
rect 13854 6025 13980 6178
rect 14046 6025 14172 6178
rect 14624 6025 14656 6178
rect 14722 6025 14848 6178
rect 14914 6025 15040 6178
rect 15106 6025 15232 6178
rect 15298 6025 15424 6178
rect 15490 6025 15616 6178
rect 15682 6025 15808 6178
rect 15874 6025 16000 6178
rect 16452 6025 16484 6178
rect 16550 6025 16676 6178
rect 16742 6025 16868 6178
rect 16934 6025 17060 6178
rect 17126 6025 17252 6178
rect 17318 6025 17444 6178
rect 17510 6025 17636 6178
rect 17702 6025 17828 6178
rect 18280 6025 18312 6178
rect 18378 6025 18504 6178
rect 18570 6025 18696 6178
rect 18762 6025 18888 6178
rect 18954 6025 19080 6178
rect 19146 6025 19272 6178
rect 19338 6025 19464 6178
rect 19530 6025 19656 6178
rect 20108 6025 20140 6178
rect 20206 6025 20332 6178
rect 20398 6025 20524 6178
rect 20590 6025 20716 6178
rect 20782 6025 20908 6178
rect 20974 6025 21100 6178
rect 21166 6025 21292 6178
rect 21358 6025 21484 6178
rect 32 6015 98 6025
rect 224 6015 290 6025
rect 416 6015 482 6025
rect 608 6015 674 6025
rect 800 6015 866 6025
rect 992 6015 1058 6025
rect 1184 6015 1250 6025
rect 1376 6015 1442 6025
rect 1860 6015 1926 6025
rect 2052 6015 2118 6025
rect 2244 6015 2310 6025
rect 2436 6015 2502 6025
rect 2628 6015 2694 6025
rect 2820 6015 2886 6025
rect 3012 6015 3078 6025
rect 3204 6015 3270 6025
rect 3688 6015 3754 6025
rect 3880 6015 3946 6025
rect 4072 6015 4138 6025
rect 4264 6015 4330 6025
rect 4456 6015 4522 6025
rect 4648 6015 4714 6025
rect 4840 6015 4906 6025
rect 5032 6015 5098 6025
rect 5516 6015 5582 6025
rect 5708 6015 5774 6025
rect 5900 6015 5966 6025
rect 6092 6015 6158 6025
rect 6284 6015 6350 6025
rect 6476 6015 6542 6025
rect 6668 6015 6734 6025
rect 6860 6015 6926 6025
rect 7344 6015 7410 6025
rect 7536 6015 7602 6025
rect 7728 6015 7794 6025
rect 7920 6015 7986 6025
rect 8112 6015 8178 6025
rect 8304 6015 8370 6025
rect 8496 6015 8562 6025
rect 8688 6015 8754 6025
rect 9172 6015 9238 6025
rect 9364 6015 9430 6025
rect 9556 6015 9622 6025
rect 9748 6015 9814 6025
rect 9940 6015 10006 6025
rect 10132 6015 10198 6025
rect 10324 6015 10390 6025
rect 10516 6015 10582 6025
rect 11000 6015 11066 6025
rect 11192 6015 11258 6025
rect 11384 6015 11450 6025
rect 11576 6015 11642 6025
rect 11768 6015 11834 6025
rect 11960 6015 12026 6025
rect 12152 6015 12218 6025
rect 12344 6015 12410 6025
rect 12828 6015 12894 6025
rect 13020 6015 13086 6025
rect 13212 6015 13278 6025
rect 13404 6015 13470 6025
rect 13596 6015 13662 6025
rect 13788 6015 13854 6025
rect 13980 6015 14046 6025
rect 14172 6015 14238 6025
rect 14656 6015 14722 6025
rect 14848 6015 14914 6025
rect 15040 6015 15106 6025
rect 15232 6015 15298 6025
rect 15424 6015 15490 6025
rect 15616 6015 15682 6025
rect 15808 6015 15874 6025
rect 16000 6015 16066 6025
rect 16484 6015 16550 6025
rect 16676 6015 16742 6025
rect 16868 6015 16934 6025
rect 17060 6015 17126 6025
rect 17252 6015 17318 6025
rect 17444 6015 17510 6025
rect 17636 6015 17702 6025
rect 17828 6015 17894 6025
rect 18312 6015 18378 6025
rect 18504 6015 18570 6025
rect 18696 6015 18762 6025
rect 18888 6015 18954 6025
rect 19080 6015 19146 6025
rect 19272 6015 19338 6025
rect 19464 6015 19530 6025
rect 19656 6015 19722 6025
rect 20140 6015 20206 6025
rect 20332 6015 20398 6025
rect 20524 6015 20590 6025
rect 20716 6015 20782 6025
rect 20908 6015 20974 6025
rect 21100 6015 21166 6025
rect 21292 6015 21358 6025
rect 21484 6015 21550 6025
rect 128 5965 194 5975
rect 320 5965 386 5975
rect 512 5965 578 5975
rect 704 5965 770 5975
rect 896 5965 962 5975
rect 1088 5965 1154 5975
rect 1280 5965 1346 5975
rect 1472 5965 1528 5975
rect 1956 5965 2022 5975
rect 2148 5965 2214 5975
rect 2340 5965 2406 5975
rect 2532 5965 2598 5975
rect 2724 5965 2790 5975
rect 2916 5965 2982 5975
rect 3108 5965 3174 5975
rect 3300 5965 3356 5975
rect 3784 5965 3850 5975
rect 3976 5965 4042 5975
rect 4168 5965 4234 5975
rect 4360 5965 4426 5975
rect 4552 5965 4618 5975
rect 4744 5965 4810 5975
rect 4936 5965 5002 5975
rect 5128 5965 5184 5975
rect 5612 5965 5678 5975
rect 5804 5965 5870 5975
rect 5996 5965 6062 5975
rect 6188 5965 6254 5975
rect 6380 5965 6446 5975
rect 6572 5965 6638 5975
rect 6764 5965 6830 5975
rect 6956 5965 7012 5975
rect 7440 5965 7506 5975
rect 7632 5965 7698 5975
rect 7824 5965 7890 5975
rect 8016 5965 8082 5975
rect 8208 5965 8274 5975
rect 8400 5965 8466 5975
rect 8592 5965 8658 5975
rect 8784 5965 8840 5975
rect 9268 5965 9334 5975
rect 9460 5965 9526 5975
rect 9652 5965 9718 5975
rect 9844 5965 9910 5975
rect 10036 5965 10102 5975
rect 10228 5965 10294 5975
rect 10420 5965 10486 5975
rect 10612 5965 10668 5975
rect 11096 5965 11162 5975
rect 11288 5965 11354 5975
rect 11480 5965 11546 5975
rect 11672 5965 11738 5975
rect 11864 5965 11930 5975
rect 12056 5965 12122 5975
rect 12248 5965 12314 5975
rect 12440 5965 12496 5975
rect 12924 5965 12990 5975
rect 13116 5965 13182 5975
rect 13308 5965 13374 5975
rect 13500 5965 13566 5975
rect 13692 5965 13758 5975
rect 13884 5965 13950 5975
rect 14076 5965 14142 5975
rect 14268 5965 14324 5975
rect 14752 5965 14818 5975
rect 14944 5965 15010 5975
rect 15136 5965 15202 5975
rect 15328 5965 15394 5975
rect 15520 5965 15586 5975
rect 15712 5965 15778 5975
rect 15904 5965 15970 5975
rect 16096 5965 16152 5975
rect 16580 5965 16646 5975
rect 16772 5965 16838 5975
rect 16964 5965 17030 5975
rect 17156 5965 17222 5975
rect 17348 5965 17414 5975
rect 17540 5965 17606 5975
rect 17732 5965 17798 5975
rect 17924 5965 17980 5975
rect 18408 5965 18474 5975
rect 18600 5965 18666 5975
rect 18792 5965 18858 5975
rect 18984 5965 19050 5975
rect 19176 5965 19242 5975
rect 19368 5965 19434 5975
rect 19560 5965 19626 5975
rect 19752 5965 19808 5975
rect 20236 5965 20302 5975
rect 20428 5965 20494 5975
rect 20620 5965 20686 5975
rect 20812 5965 20878 5975
rect 21004 5965 21070 5975
rect 21196 5965 21262 5975
rect 21388 5965 21454 5975
rect 21580 5965 21636 5975
rect 0 5812 128 5965
rect 194 5812 320 5965
rect 386 5812 512 5965
rect 578 5812 704 5965
rect 770 5812 896 5965
rect 962 5812 1088 5965
rect 1154 5812 1280 5965
rect 1346 5812 1472 5965
rect 1528 5812 1708 5965
rect 1828 5812 1956 5965
rect 2022 5812 2148 5965
rect 2214 5812 2340 5965
rect 2406 5812 2532 5965
rect 2598 5812 2724 5965
rect 2790 5812 2916 5965
rect 2982 5812 3108 5965
rect 3174 5812 3300 5965
rect 3356 5812 3536 5965
rect 3656 5812 3784 5965
rect 3850 5812 3976 5965
rect 4042 5812 4168 5965
rect 4234 5812 4360 5965
rect 4426 5812 4552 5965
rect 4618 5812 4744 5965
rect 4810 5812 4936 5965
rect 5002 5812 5128 5965
rect 5184 5812 5364 5965
rect 5484 5812 5612 5965
rect 5678 5812 5804 5965
rect 5870 5812 5996 5965
rect 6062 5812 6188 5965
rect 6254 5812 6380 5965
rect 6446 5812 6572 5965
rect 6638 5812 6764 5965
rect 6830 5812 6956 5965
rect 7012 5812 7192 5965
rect 7312 5812 7440 5965
rect 7506 5812 7632 5965
rect 7698 5812 7824 5965
rect 7890 5812 8016 5965
rect 8082 5812 8208 5965
rect 8274 5812 8400 5965
rect 8466 5812 8592 5965
rect 8658 5812 8784 5965
rect 8840 5812 9020 5965
rect 9140 5812 9268 5965
rect 9334 5812 9460 5965
rect 9526 5812 9652 5965
rect 9718 5812 9844 5965
rect 9910 5812 10036 5965
rect 10102 5812 10228 5965
rect 10294 5812 10420 5965
rect 10486 5812 10612 5965
rect 10668 5812 10848 5965
rect 10968 5812 11096 5965
rect 11162 5812 11288 5965
rect 11354 5812 11480 5965
rect 11546 5812 11672 5965
rect 11738 5812 11864 5965
rect 11930 5812 12056 5965
rect 12122 5812 12248 5965
rect 12314 5812 12440 5965
rect 12496 5812 12676 5965
rect 12796 5812 12924 5965
rect 12990 5812 13116 5965
rect 13182 5812 13308 5965
rect 13374 5812 13500 5965
rect 13566 5812 13692 5965
rect 13758 5812 13884 5965
rect 13950 5812 14076 5965
rect 14142 5812 14268 5965
rect 14324 5812 14504 5965
rect 14624 5812 14752 5965
rect 14818 5812 14944 5965
rect 15010 5812 15136 5965
rect 15202 5812 15328 5965
rect 15394 5812 15520 5965
rect 15586 5812 15712 5965
rect 15778 5812 15904 5965
rect 15970 5812 16096 5965
rect 16152 5812 16332 5965
rect 16452 5812 16580 5965
rect 16646 5812 16772 5965
rect 16838 5812 16964 5965
rect 17030 5812 17156 5965
rect 17222 5812 17348 5965
rect 17414 5812 17540 5965
rect 17606 5812 17732 5965
rect 17798 5812 17924 5965
rect 17980 5812 18160 5965
rect 18280 5812 18408 5965
rect 18474 5812 18600 5965
rect 18666 5812 18792 5965
rect 18858 5812 18984 5965
rect 19050 5812 19176 5965
rect 19242 5812 19368 5965
rect 19434 5812 19560 5965
rect 19626 5812 19752 5965
rect 19808 5812 19988 5965
rect 20108 5812 20236 5965
rect 20302 5812 20428 5965
rect 20494 5812 20620 5965
rect 20686 5812 20812 5965
rect 20878 5812 21004 5965
rect 21070 5812 21196 5965
rect 21262 5812 21388 5965
rect 21454 5812 21580 5965
rect 21636 5812 21816 5965
rect 128 5802 194 5812
rect 320 5802 386 5812
rect 512 5802 578 5812
rect 704 5802 770 5812
rect 896 5802 962 5812
rect 1088 5802 1154 5812
rect 1280 5802 1346 5812
rect 1472 5802 1528 5812
rect 1956 5802 2022 5812
rect 2148 5802 2214 5812
rect 2340 5802 2406 5812
rect 2532 5802 2598 5812
rect 2724 5802 2790 5812
rect 2916 5802 2982 5812
rect 3108 5802 3174 5812
rect 3300 5802 3356 5812
rect 3784 5802 3850 5812
rect 3976 5802 4042 5812
rect 4168 5802 4234 5812
rect 4360 5802 4426 5812
rect 4552 5802 4618 5812
rect 4744 5802 4810 5812
rect 4936 5802 5002 5812
rect 5128 5802 5184 5812
rect 5612 5802 5678 5812
rect 5804 5802 5870 5812
rect 5996 5802 6062 5812
rect 6188 5802 6254 5812
rect 6380 5802 6446 5812
rect 6572 5802 6638 5812
rect 6764 5802 6830 5812
rect 6956 5802 7012 5812
rect 7440 5802 7506 5812
rect 7632 5802 7698 5812
rect 7824 5802 7890 5812
rect 8016 5802 8082 5812
rect 8208 5802 8274 5812
rect 8400 5802 8466 5812
rect 8592 5802 8658 5812
rect 8784 5802 8840 5812
rect 9268 5802 9334 5812
rect 9460 5802 9526 5812
rect 9652 5802 9718 5812
rect 9844 5802 9910 5812
rect 10036 5802 10102 5812
rect 10228 5802 10294 5812
rect 10420 5802 10486 5812
rect 10612 5802 10668 5812
rect 11096 5802 11162 5812
rect 11288 5802 11354 5812
rect 11480 5802 11546 5812
rect 11672 5802 11738 5812
rect 11864 5802 11930 5812
rect 12056 5802 12122 5812
rect 12248 5802 12314 5812
rect 12440 5802 12496 5812
rect 12924 5802 12990 5812
rect 13116 5802 13182 5812
rect 13308 5802 13374 5812
rect 13500 5802 13566 5812
rect 13692 5802 13758 5812
rect 13884 5802 13950 5812
rect 14076 5802 14142 5812
rect 14268 5802 14324 5812
rect 14752 5802 14818 5812
rect 14944 5802 15010 5812
rect 15136 5802 15202 5812
rect 15328 5802 15394 5812
rect 15520 5802 15586 5812
rect 15712 5802 15778 5812
rect 15904 5802 15970 5812
rect 16096 5802 16152 5812
rect 16580 5802 16646 5812
rect 16772 5802 16838 5812
rect 16964 5802 17030 5812
rect 17156 5802 17222 5812
rect 17348 5802 17414 5812
rect 17540 5802 17606 5812
rect 17732 5802 17798 5812
rect 17924 5802 17980 5812
rect 18408 5802 18474 5812
rect 18600 5802 18666 5812
rect 18792 5802 18858 5812
rect 18984 5802 19050 5812
rect 19176 5802 19242 5812
rect 19368 5802 19434 5812
rect 19560 5802 19626 5812
rect 19752 5802 19808 5812
rect 20236 5802 20302 5812
rect 20428 5802 20494 5812
rect 20620 5802 20686 5812
rect 20812 5802 20878 5812
rect 21004 5802 21070 5812
rect 21196 5802 21262 5812
rect 21388 5802 21454 5812
rect 21580 5802 21636 5812
rect 32 5464 98 5474
rect 224 5464 290 5474
rect 416 5464 482 5474
rect 608 5464 674 5474
rect 800 5464 866 5474
rect 992 5464 1058 5474
rect 1184 5464 1250 5474
rect 1376 5464 1442 5474
rect 1860 5464 1926 5474
rect 2052 5464 2118 5474
rect 2244 5464 2310 5474
rect 2436 5464 2502 5474
rect 2628 5464 2694 5474
rect 2820 5464 2886 5474
rect 3012 5464 3078 5474
rect 3204 5464 3270 5474
rect 3688 5464 3754 5474
rect 3880 5464 3946 5474
rect 4072 5464 4138 5474
rect 4264 5464 4330 5474
rect 4456 5464 4522 5474
rect 4648 5464 4714 5474
rect 4840 5464 4906 5474
rect 5032 5464 5098 5474
rect 5516 5464 5582 5474
rect 5708 5464 5774 5474
rect 5900 5464 5966 5474
rect 6092 5464 6158 5474
rect 6284 5464 6350 5474
rect 6476 5464 6542 5474
rect 6668 5464 6734 5474
rect 6860 5464 6926 5474
rect 7344 5464 7410 5474
rect 7536 5464 7602 5474
rect 7728 5464 7794 5474
rect 7920 5464 7986 5474
rect 8112 5464 8178 5474
rect 8304 5464 8370 5474
rect 8496 5464 8562 5474
rect 8688 5464 8754 5474
rect 9172 5464 9238 5474
rect 9364 5464 9430 5474
rect 9556 5464 9622 5474
rect 9748 5464 9814 5474
rect 9940 5464 10006 5474
rect 10132 5464 10198 5474
rect 10324 5464 10390 5474
rect 10516 5464 10582 5474
rect 11000 5464 11066 5474
rect 11192 5464 11258 5474
rect 11384 5464 11450 5474
rect 11576 5464 11642 5474
rect 11768 5464 11834 5474
rect 11960 5464 12026 5474
rect 12152 5464 12218 5474
rect 12344 5464 12410 5474
rect 12828 5464 12894 5474
rect 13020 5464 13086 5474
rect 13212 5464 13278 5474
rect 13404 5464 13470 5474
rect 13596 5464 13662 5474
rect 13788 5464 13854 5474
rect 13980 5464 14046 5474
rect 14172 5464 14238 5474
rect 14656 5464 14722 5474
rect 14848 5464 14914 5474
rect 15040 5464 15106 5474
rect 15232 5464 15298 5474
rect 15424 5464 15490 5474
rect 15616 5464 15682 5474
rect 15808 5464 15874 5474
rect 16000 5464 16066 5474
rect 16484 5464 16550 5474
rect 16676 5464 16742 5474
rect 16868 5464 16934 5474
rect 17060 5464 17126 5474
rect 17252 5464 17318 5474
rect 17444 5464 17510 5474
rect 17636 5464 17702 5474
rect 17828 5464 17894 5474
rect 18312 5464 18378 5474
rect 18504 5464 18570 5474
rect 18696 5464 18762 5474
rect 18888 5464 18954 5474
rect 19080 5464 19146 5474
rect 19272 5464 19338 5474
rect 19464 5464 19530 5474
rect 19656 5464 19722 5474
rect 20140 5464 20206 5474
rect 20332 5464 20398 5474
rect 20524 5464 20590 5474
rect 20716 5464 20782 5474
rect 20908 5464 20974 5474
rect 21100 5464 21166 5474
rect 21292 5464 21358 5474
rect 21484 5464 21550 5474
rect 0 5311 32 5464
rect 98 5311 224 5464
rect 290 5311 416 5464
rect 482 5311 608 5464
rect 674 5311 800 5464
rect 866 5311 992 5464
rect 1058 5311 1184 5464
rect 1250 5311 1376 5464
rect 1828 5311 1860 5464
rect 1926 5311 2052 5464
rect 2118 5311 2244 5464
rect 2310 5311 2436 5464
rect 2502 5311 2628 5464
rect 2694 5311 2820 5464
rect 2886 5311 3012 5464
rect 3078 5311 3204 5464
rect 3656 5311 3688 5464
rect 3754 5311 3880 5464
rect 3946 5311 4072 5464
rect 4138 5311 4264 5464
rect 4330 5311 4456 5464
rect 4522 5311 4648 5464
rect 4714 5311 4840 5464
rect 4906 5311 5032 5464
rect 5484 5311 5516 5464
rect 5582 5311 5708 5464
rect 5774 5311 5900 5464
rect 5966 5311 6092 5464
rect 6158 5311 6284 5464
rect 6350 5311 6476 5464
rect 6542 5311 6668 5464
rect 6734 5311 6860 5464
rect 7312 5311 7344 5464
rect 7410 5311 7536 5464
rect 7602 5311 7728 5464
rect 7794 5311 7920 5464
rect 7986 5311 8112 5464
rect 8178 5311 8304 5464
rect 8370 5311 8496 5464
rect 8562 5311 8688 5464
rect 9140 5311 9172 5464
rect 9238 5311 9364 5464
rect 9430 5311 9556 5464
rect 9622 5311 9748 5464
rect 9814 5311 9940 5464
rect 10006 5311 10132 5464
rect 10198 5311 10324 5464
rect 10390 5311 10516 5464
rect 10968 5311 11000 5464
rect 11066 5311 11192 5464
rect 11258 5311 11384 5464
rect 11450 5311 11576 5464
rect 11642 5311 11768 5464
rect 11834 5311 11960 5464
rect 12026 5311 12152 5464
rect 12218 5311 12344 5464
rect 12796 5311 12828 5464
rect 12894 5311 13020 5464
rect 13086 5311 13212 5464
rect 13278 5311 13404 5464
rect 13470 5311 13596 5464
rect 13662 5311 13788 5464
rect 13854 5311 13980 5464
rect 14046 5311 14172 5464
rect 14624 5311 14656 5464
rect 14722 5311 14848 5464
rect 14914 5311 15040 5464
rect 15106 5311 15232 5464
rect 15298 5311 15424 5464
rect 15490 5311 15616 5464
rect 15682 5311 15808 5464
rect 15874 5311 16000 5464
rect 16452 5311 16484 5464
rect 16550 5311 16676 5464
rect 16742 5311 16868 5464
rect 16934 5311 17060 5464
rect 17126 5311 17252 5464
rect 17318 5311 17444 5464
rect 17510 5311 17636 5464
rect 17702 5311 17828 5464
rect 18280 5311 18312 5464
rect 18378 5311 18504 5464
rect 18570 5311 18696 5464
rect 18762 5311 18888 5464
rect 18954 5311 19080 5464
rect 19146 5311 19272 5464
rect 19338 5311 19464 5464
rect 19530 5311 19656 5464
rect 20108 5311 20140 5464
rect 20206 5311 20332 5464
rect 20398 5311 20524 5464
rect 20590 5311 20716 5464
rect 20782 5311 20908 5464
rect 20974 5311 21100 5464
rect 21166 5311 21292 5464
rect 21358 5311 21484 5464
rect 32 5301 98 5311
rect 224 5301 290 5311
rect 416 5301 482 5311
rect 608 5301 674 5311
rect 800 5301 866 5311
rect 992 5301 1058 5311
rect 1184 5301 1250 5311
rect 1376 5301 1442 5311
rect 1860 5301 1926 5311
rect 2052 5301 2118 5311
rect 2244 5301 2310 5311
rect 2436 5301 2502 5311
rect 2628 5301 2694 5311
rect 2820 5301 2886 5311
rect 3012 5301 3078 5311
rect 3204 5301 3270 5311
rect 3688 5301 3754 5311
rect 3880 5301 3946 5311
rect 4072 5301 4138 5311
rect 4264 5301 4330 5311
rect 4456 5301 4522 5311
rect 4648 5301 4714 5311
rect 4840 5301 4906 5311
rect 5032 5301 5098 5311
rect 5516 5301 5582 5311
rect 5708 5301 5774 5311
rect 5900 5301 5966 5311
rect 6092 5301 6158 5311
rect 6284 5301 6350 5311
rect 6476 5301 6542 5311
rect 6668 5301 6734 5311
rect 6860 5301 6926 5311
rect 7344 5301 7410 5311
rect 7536 5301 7602 5311
rect 7728 5301 7794 5311
rect 7920 5301 7986 5311
rect 8112 5301 8178 5311
rect 8304 5301 8370 5311
rect 8496 5301 8562 5311
rect 8688 5301 8754 5311
rect 9172 5301 9238 5311
rect 9364 5301 9430 5311
rect 9556 5301 9622 5311
rect 9748 5301 9814 5311
rect 9940 5301 10006 5311
rect 10132 5301 10198 5311
rect 10324 5301 10390 5311
rect 10516 5301 10582 5311
rect 11000 5301 11066 5311
rect 11192 5301 11258 5311
rect 11384 5301 11450 5311
rect 11576 5301 11642 5311
rect 11768 5301 11834 5311
rect 11960 5301 12026 5311
rect 12152 5301 12218 5311
rect 12344 5301 12410 5311
rect 12828 5301 12894 5311
rect 13020 5301 13086 5311
rect 13212 5301 13278 5311
rect 13404 5301 13470 5311
rect 13596 5301 13662 5311
rect 13788 5301 13854 5311
rect 13980 5301 14046 5311
rect 14172 5301 14238 5311
rect 14656 5301 14722 5311
rect 14848 5301 14914 5311
rect 15040 5301 15106 5311
rect 15232 5301 15298 5311
rect 15424 5301 15490 5311
rect 15616 5301 15682 5311
rect 15808 5301 15874 5311
rect 16000 5301 16066 5311
rect 16484 5301 16550 5311
rect 16676 5301 16742 5311
rect 16868 5301 16934 5311
rect 17060 5301 17126 5311
rect 17252 5301 17318 5311
rect 17444 5301 17510 5311
rect 17636 5301 17702 5311
rect 17828 5301 17894 5311
rect 18312 5301 18378 5311
rect 18504 5301 18570 5311
rect 18696 5301 18762 5311
rect 18888 5301 18954 5311
rect 19080 5301 19146 5311
rect 19272 5301 19338 5311
rect 19464 5301 19530 5311
rect 19656 5301 19722 5311
rect 20140 5301 20206 5311
rect 20332 5301 20398 5311
rect 20524 5301 20590 5311
rect 20716 5301 20782 5311
rect 20908 5301 20974 5311
rect 21100 5301 21166 5311
rect 21292 5301 21358 5311
rect 21484 5301 21550 5311
rect 128 5251 194 5261
rect 320 5251 386 5261
rect 512 5251 578 5261
rect 704 5251 770 5261
rect 896 5251 962 5261
rect 1088 5251 1154 5261
rect 1280 5251 1346 5261
rect 1472 5251 1528 5261
rect 1956 5251 2022 5261
rect 2148 5251 2214 5261
rect 2340 5251 2406 5261
rect 2532 5251 2598 5261
rect 2724 5251 2790 5261
rect 2916 5251 2982 5261
rect 3108 5251 3174 5261
rect 3300 5251 3356 5261
rect 3784 5251 3850 5261
rect 3976 5251 4042 5261
rect 4168 5251 4234 5261
rect 4360 5251 4426 5261
rect 4552 5251 4618 5261
rect 4744 5251 4810 5261
rect 4936 5251 5002 5261
rect 5128 5251 5184 5261
rect 5612 5251 5678 5261
rect 5804 5251 5870 5261
rect 5996 5251 6062 5261
rect 6188 5251 6254 5261
rect 6380 5251 6446 5261
rect 6572 5251 6638 5261
rect 6764 5251 6830 5261
rect 6956 5251 7012 5261
rect 7440 5251 7506 5261
rect 7632 5251 7698 5261
rect 7824 5251 7890 5261
rect 8016 5251 8082 5261
rect 8208 5251 8274 5261
rect 8400 5251 8466 5261
rect 8592 5251 8658 5261
rect 8784 5251 8840 5261
rect 9268 5251 9334 5261
rect 9460 5251 9526 5261
rect 9652 5251 9718 5261
rect 9844 5251 9910 5261
rect 10036 5251 10102 5261
rect 10228 5251 10294 5261
rect 10420 5251 10486 5261
rect 10612 5251 10668 5261
rect 11096 5251 11162 5261
rect 11288 5251 11354 5261
rect 11480 5251 11546 5261
rect 11672 5251 11738 5261
rect 11864 5251 11930 5261
rect 12056 5251 12122 5261
rect 12248 5251 12314 5261
rect 12440 5251 12496 5261
rect 12924 5251 12990 5261
rect 13116 5251 13182 5261
rect 13308 5251 13374 5261
rect 13500 5251 13566 5261
rect 13692 5251 13758 5261
rect 13884 5251 13950 5261
rect 14076 5251 14142 5261
rect 14268 5251 14324 5261
rect 14752 5251 14818 5261
rect 14944 5251 15010 5261
rect 15136 5251 15202 5261
rect 15328 5251 15394 5261
rect 15520 5251 15586 5261
rect 15712 5251 15778 5261
rect 15904 5251 15970 5261
rect 16096 5251 16152 5261
rect 16580 5251 16646 5261
rect 16772 5251 16838 5261
rect 16964 5251 17030 5261
rect 17156 5251 17222 5261
rect 17348 5251 17414 5261
rect 17540 5251 17606 5261
rect 17732 5251 17798 5261
rect 17924 5251 17980 5261
rect 18408 5251 18474 5261
rect 18600 5251 18666 5261
rect 18792 5251 18858 5261
rect 18984 5251 19050 5261
rect 19176 5251 19242 5261
rect 19368 5251 19434 5261
rect 19560 5251 19626 5261
rect 19752 5251 19808 5261
rect 20236 5251 20302 5261
rect 20428 5251 20494 5261
rect 20620 5251 20686 5261
rect 20812 5251 20878 5261
rect 21004 5251 21070 5261
rect 21196 5251 21262 5261
rect 21388 5251 21454 5261
rect 21580 5251 21636 5261
rect 0 5098 128 5251
rect 194 5098 320 5251
rect 386 5098 512 5251
rect 578 5098 704 5251
rect 770 5098 896 5251
rect 962 5098 1088 5251
rect 1154 5098 1280 5251
rect 1346 5098 1472 5251
rect 1528 5098 1708 5251
rect 1828 5098 1956 5251
rect 2022 5098 2148 5251
rect 2214 5098 2340 5251
rect 2406 5098 2532 5251
rect 2598 5098 2724 5251
rect 2790 5098 2916 5251
rect 2982 5098 3108 5251
rect 3174 5098 3300 5251
rect 3356 5098 3536 5251
rect 3656 5098 3784 5251
rect 3850 5098 3976 5251
rect 4042 5098 4168 5251
rect 4234 5098 4360 5251
rect 4426 5098 4552 5251
rect 4618 5098 4744 5251
rect 4810 5098 4936 5251
rect 5002 5098 5128 5251
rect 5184 5098 5364 5251
rect 5484 5098 5612 5251
rect 5678 5098 5804 5251
rect 5870 5098 5996 5251
rect 6062 5098 6188 5251
rect 6254 5098 6380 5251
rect 6446 5098 6572 5251
rect 6638 5098 6764 5251
rect 6830 5098 6956 5251
rect 7012 5098 7192 5251
rect 7312 5098 7440 5251
rect 7506 5098 7632 5251
rect 7698 5098 7824 5251
rect 7890 5098 8016 5251
rect 8082 5098 8208 5251
rect 8274 5098 8400 5251
rect 8466 5098 8592 5251
rect 8658 5098 8784 5251
rect 8840 5098 9020 5251
rect 9140 5098 9268 5251
rect 9334 5098 9460 5251
rect 9526 5098 9652 5251
rect 9718 5098 9844 5251
rect 9910 5098 10036 5251
rect 10102 5098 10228 5251
rect 10294 5098 10420 5251
rect 10486 5098 10612 5251
rect 10668 5098 10848 5251
rect 10968 5098 11096 5251
rect 11162 5098 11288 5251
rect 11354 5098 11480 5251
rect 11546 5098 11672 5251
rect 11738 5098 11864 5251
rect 11930 5098 12056 5251
rect 12122 5098 12248 5251
rect 12314 5098 12440 5251
rect 12496 5098 12676 5251
rect 12796 5098 12924 5251
rect 12990 5098 13116 5251
rect 13182 5098 13308 5251
rect 13374 5098 13500 5251
rect 13566 5098 13692 5251
rect 13758 5098 13884 5251
rect 13950 5098 14076 5251
rect 14142 5098 14268 5251
rect 14324 5098 14504 5251
rect 14624 5098 14752 5251
rect 14818 5098 14944 5251
rect 15010 5098 15136 5251
rect 15202 5098 15328 5251
rect 15394 5098 15520 5251
rect 15586 5098 15712 5251
rect 15778 5098 15904 5251
rect 15970 5098 16096 5251
rect 16152 5098 16332 5251
rect 16452 5098 16580 5251
rect 16646 5098 16772 5251
rect 16838 5098 16964 5251
rect 17030 5098 17156 5251
rect 17222 5098 17348 5251
rect 17414 5098 17540 5251
rect 17606 5098 17732 5251
rect 17798 5098 17924 5251
rect 17980 5098 18160 5251
rect 18280 5098 18408 5251
rect 18474 5098 18600 5251
rect 18666 5098 18792 5251
rect 18858 5098 18984 5251
rect 19050 5098 19176 5251
rect 19242 5098 19368 5251
rect 19434 5098 19560 5251
rect 19626 5098 19752 5251
rect 19808 5098 19988 5251
rect 20108 5098 20236 5251
rect 20302 5098 20428 5251
rect 20494 5098 20620 5251
rect 20686 5098 20812 5251
rect 20878 5098 21004 5251
rect 21070 5098 21196 5251
rect 21262 5098 21388 5251
rect 21454 5098 21580 5251
rect 21636 5098 21816 5251
rect 128 5088 194 5098
rect 320 5088 386 5098
rect 512 5088 578 5098
rect 704 5088 770 5098
rect 896 5088 962 5098
rect 1088 5088 1154 5098
rect 1280 5088 1346 5098
rect 1472 5088 1528 5098
rect 1956 5088 2022 5098
rect 2148 5088 2214 5098
rect 2340 5088 2406 5098
rect 2532 5088 2598 5098
rect 2724 5088 2790 5098
rect 2916 5088 2982 5098
rect 3108 5088 3174 5098
rect 3300 5088 3356 5098
rect 3784 5088 3850 5098
rect 3976 5088 4042 5098
rect 4168 5088 4234 5098
rect 4360 5088 4426 5098
rect 4552 5088 4618 5098
rect 4744 5088 4810 5098
rect 4936 5088 5002 5098
rect 5128 5088 5184 5098
rect 5612 5088 5678 5098
rect 5804 5088 5870 5098
rect 5996 5088 6062 5098
rect 6188 5088 6254 5098
rect 6380 5088 6446 5098
rect 6572 5088 6638 5098
rect 6764 5088 6830 5098
rect 6956 5088 7012 5098
rect 7440 5088 7506 5098
rect 7632 5088 7698 5098
rect 7824 5088 7890 5098
rect 8016 5088 8082 5098
rect 8208 5088 8274 5098
rect 8400 5088 8466 5098
rect 8592 5088 8658 5098
rect 8784 5088 8840 5098
rect 9268 5088 9334 5098
rect 9460 5088 9526 5098
rect 9652 5088 9718 5098
rect 9844 5088 9910 5098
rect 10036 5088 10102 5098
rect 10228 5088 10294 5098
rect 10420 5088 10486 5098
rect 10612 5088 10668 5098
rect 11096 5088 11162 5098
rect 11288 5088 11354 5098
rect 11480 5088 11546 5098
rect 11672 5088 11738 5098
rect 11864 5088 11930 5098
rect 12056 5088 12122 5098
rect 12248 5088 12314 5098
rect 12440 5088 12496 5098
rect 12924 5088 12990 5098
rect 13116 5088 13182 5098
rect 13308 5088 13374 5098
rect 13500 5088 13566 5098
rect 13692 5088 13758 5098
rect 13884 5088 13950 5098
rect 14076 5088 14142 5098
rect 14268 5088 14324 5098
rect 14752 5088 14818 5098
rect 14944 5088 15010 5098
rect 15136 5088 15202 5098
rect 15328 5088 15394 5098
rect 15520 5088 15586 5098
rect 15712 5088 15778 5098
rect 15904 5088 15970 5098
rect 16096 5088 16152 5098
rect 16580 5088 16646 5098
rect 16772 5088 16838 5098
rect 16964 5088 17030 5098
rect 17156 5088 17222 5098
rect 17348 5088 17414 5098
rect 17540 5088 17606 5098
rect 17732 5088 17798 5098
rect 17924 5088 17980 5098
rect 18408 5088 18474 5098
rect 18600 5088 18666 5098
rect 18792 5088 18858 5098
rect 18984 5088 19050 5098
rect 19176 5088 19242 5098
rect 19368 5088 19434 5098
rect 19560 5088 19626 5098
rect 19752 5088 19808 5098
rect 20236 5088 20302 5098
rect 20428 5088 20494 5098
rect 20620 5088 20686 5098
rect 20812 5088 20878 5098
rect 21004 5088 21070 5098
rect 21196 5088 21262 5098
rect 21388 5088 21454 5098
rect 21580 5088 21636 5098
rect 32 4750 98 4760
rect 224 4750 290 4760
rect 416 4750 482 4760
rect 608 4750 674 4760
rect 800 4750 866 4760
rect 992 4750 1058 4760
rect 1184 4750 1250 4760
rect 1376 4750 1442 4760
rect 1860 4750 1926 4760
rect 2052 4750 2118 4760
rect 2244 4750 2310 4760
rect 2436 4750 2502 4760
rect 2628 4750 2694 4760
rect 2820 4750 2886 4760
rect 3012 4750 3078 4760
rect 3204 4750 3270 4760
rect 3688 4750 3754 4760
rect 3880 4750 3946 4760
rect 4072 4750 4138 4760
rect 4264 4750 4330 4760
rect 4456 4750 4522 4760
rect 4648 4750 4714 4760
rect 4840 4750 4906 4760
rect 5032 4750 5098 4760
rect 5516 4750 5582 4760
rect 5708 4750 5774 4760
rect 5900 4750 5966 4760
rect 6092 4750 6158 4760
rect 6284 4750 6350 4760
rect 6476 4750 6542 4760
rect 6668 4750 6734 4760
rect 6860 4750 6926 4760
rect 7344 4750 7410 4760
rect 7536 4750 7602 4760
rect 7728 4750 7794 4760
rect 7920 4750 7986 4760
rect 8112 4750 8178 4760
rect 8304 4750 8370 4760
rect 8496 4750 8562 4760
rect 8688 4750 8754 4760
rect 9172 4750 9238 4760
rect 9364 4750 9430 4760
rect 9556 4750 9622 4760
rect 9748 4750 9814 4760
rect 9940 4750 10006 4760
rect 10132 4750 10198 4760
rect 10324 4750 10390 4760
rect 10516 4750 10582 4760
rect 11000 4750 11066 4760
rect 11192 4750 11258 4760
rect 11384 4750 11450 4760
rect 11576 4750 11642 4760
rect 11768 4750 11834 4760
rect 11960 4750 12026 4760
rect 12152 4750 12218 4760
rect 12344 4750 12410 4760
rect 12828 4750 12894 4760
rect 13020 4750 13086 4760
rect 13212 4750 13278 4760
rect 13404 4750 13470 4760
rect 13596 4750 13662 4760
rect 13788 4750 13854 4760
rect 13980 4750 14046 4760
rect 14172 4750 14238 4760
rect 14656 4750 14722 4760
rect 14848 4750 14914 4760
rect 15040 4750 15106 4760
rect 15232 4750 15298 4760
rect 15424 4750 15490 4760
rect 15616 4750 15682 4760
rect 15808 4750 15874 4760
rect 16000 4750 16066 4760
rect 16484 4750 16550 4760
rect 16676 4750 16742 4760
rect 16868 4750 16934 4760
rect 17060 4750 17126 4760
rect 17252 4750 17318 4760
rect 17444 4750 17510 4760
rect 17636 4750 17702 4760
rect 17828 4750 17894 4760
rect 18312 4750 18378 4760
rect 18504 4750 18570 4760
rect 18696 4750 18762 4760
rect 18888 4750 18954 4760
rect 19080 4750 19146 4760
rect 19272 4750 19338 4760
rect 19464 4750 19530 4760
rect 19656 4750 19722 4760
rect 20140 4750 20206 4760
rect 20332 4750 20398 4760
rect 20524 4750 20590 4760
rect 20716 4750 20782 4760
rect 20908 4750 20974 4760
rect 21100 4750 21166 4760
rect 21292 4750 21358 4760
rect 21484 4750 21550 4760
rect 0 4597 32 4750
rect 98 4597 224 4750
rect 290 4597 416 4750
rect 482 4597 608 4750
rect 674 4597 800 4750
rect 866 4597 992 4750
rect 1058 4597 1184 4750
rect 1250 4597 1376 4750
rect 1828 4597 1860 4750
rect 1926 4597 2052 4750
rect 2118 4597 2244 4750
rect 2310 4597 2436 4750
rect 2502 4597 2628 4750
rect 2694 4597 2820 4750
rect 2886 4597 3012 4750
rect 3078 4597 3204 4750
rect 3656 4597 3688 4750
rect 3754 4597 3880 4750
rect 3946 4597 4072 4750
rect 4138 4597 4264 4750
rect 4330 4597 4456 4750
rect 4522 4597 4648 4750
rect 4714 4597 4840 4750
rect 4906 4597 5032 4750
rect 5484 4597 5516 4750
rect 5582 4597 5708 4750
rect 5774 4597 5900 4750
rect 5966 4597 6092 4750
rect 6158 4597 6284 4750
rect 6350 4597 6476 4750
rect 6542 4597 6668 4750
rect 6734 4597 6860 4750
rect 7312 4597 7344 4750
rect 7410 4597 7536 4750
rect 7602 4597 7728 4750
rect 7794 4597 7920 4750
rect 7986 4597 8112 4750
rect 8178 4597 8304 4750
rect 8370 4597 8496 4750
rect 8562 4597 8688 4750
rect 9140 4597 9172 4750
rect 9238 4597 9364 4750
rect 9430 4597 9556 4750
rect 9622 4597 9748 4750
rect 9814 4597 9940 4750
rect 10006 4597 10132 4750
rect 10198 4597 10324 4750
rect 10390 4597 10516 4750
rect 10968 4597 11000 4750
rect 11066 4597 11192 4750
rect 11258 4597 11384 4750
rect 11450 4597 11576 4750
rect 11642 4597 11768 4750
rect 11834 4597 11960 4750
rect 12026 4597 12152 4750
rect 12218 4597 12344 4750
rect 12796 4597 12828 4750
rect 12894 4597 13020 4750
rect 13086 4597 13212 4750
rect 13278 4597 13404 4750
rect 13470 4597 13596 4750
rect 13662 4597 13788 4750
rect 13854 4597 13980 4750
rect 14046 4597 14172 4750
rect 14624 4597 14656 4750
rect 14722 4597 14848 4750
rect 14914 4597 15040 4750
rect 15106 4597 15232 4750
rect 15298 4597 15424 4750
rect 15490 4597 15616 4750
rect 15682 4597 15808 4750
rect 15874 4597 16000 4750
rect 16452 4597 16484 4750
rect 16550 4597 16676 4750
rect 16742 4597 16868 4750
rect 16934 4597 17060 4750
rect 17126 4597 17252 4750
rect 17318 4597 17444 4750
rect 17510 4597 17636 4750
rect 17702 4597 17828 4750
rect 18280 4597 18312 4750
rect 18378 4597 18504 4750
rect 18570 4597 18696 4750
rect 18762 4597 18888 4750
rect 18954 4597 19080 4750
rect 19146 4597 19272 4750
rect 19338 4597 19464 4750
rect 19530 4597 19656 4750
rect 20108 4597 20140 4750
rect 20206 4597 20332 4750
rect 20398 4597 20524 4750
rect 20590 4597 20716 4750
rect 20782 4597 20908 4750
rect 20974 4597 21100 4750
rect 21166 4597 21292 4750
rect 21358 4597 21484 4750
rect 32 4587 98 4597
rect 224 4587 290 4597
rect 416 4587 482 4597
rect 608 4587 674 4597
rect 800 4587 866 4597
rect 992 4587 1058 4597
rect 1184 4587 1250 4597
rect 1376 4587 1442 4597
rect 1860 4587 1926 4597
rect 2052 4587 2118 4597
rect 2244 4587 2310 4597
rect 2436 4587 2502 4597
rect 2628 4587 2694 4597
rect 2820 4587 2886 4597
rect 3012 4587 3078 4597
rect 3204 4587 3270 4597
rect 3688 4587 3754 4597
rect 3880 4587 3946 4597
rect 4072 4587 4138 4597
rect 4264 4587 4330 4597
rect 4456 4587 4522 4597
rect 4648 4587 4714 4597
rect 4840 4587 4906 4597
rect 5032 4587 5098 4597
rect 5516 4587 5582 4597
rect 5708 4587 5774 4597
rect 5900 4587 5966 4597
rect 6092 4587 6158 4597
rect 6284 4587 6350 4597
rect 6476 4587 6542 4597
rect 6668 4587 6734 4597
rect 6860 4587 6926 4597
rect 7344 4587 7410 4597
rect 7536 4587 7602 4597
rect 7728 4587 7794 4597
rect 7920 4587 7986 4597
rect 8112 4587 8178 4597
rect 8304 4587 8370 4597
rect 8496 4587 8562 4597
rect 8688 4587 8754 4597
rect 9172 4587 9238 4597
rect 9364 4587 9430 4597
rect 9556 4587 9622 4597
rect 9748 4587 9814 4597
rect 9940 4587 10006 4597
rect 10132 4587 10198 4597
rect 10324 4587 10390 4597
rect 10516 4587 10582 4597
rect 11000 4587 11066 4597
rect 11192 4587 11258 4597
rect 11384 4587 11450 4597
rect 11576 4587 11642 4597
rect 11768 4587 11834 4597
rect 11960 4587 12026 4597
rect 12152 4587 12218 4597
rect 12344 4587 12410 4597
rect 12828 4587 12894 4597
rect 13020 4587 13086 4597
rect 13212 4587 13278 4597
rect 13404 4587 13470 4597
rect 13596 4587 13662 4597
rect 13788 4587 13854 4597
rect 13980 4587 14046 4597
rect 14172 4587 14238 4597
rect 14656 4587 14722 4597
rect 14848 4587 14914 4597
rect 15040 4587 15106 4597
rect 15232 4587 15298 4597
rect 15424 4587 15490 4597
rect 15616 4587 15682 4597
rect 15808 4587 15874 4597
rect 16000 4587 16066 4597
rect 16484 4587 16550 4597
rect 16676 4587 16742 4597
rect 16868 4587 16934 4597
rect 17060 4587 17126 4597
rect 17252 4587 17318 4597
rect 17444 4587 17510 4597
rect 17636 4587 17702 4597
rect 17828 4587 17894 4597
rect 18312 4587 18378 4597
rect 18504 4587 18570 4597
rect 18696 4587 18762 4597
rect 18888 4587 18954 4597
rect 19080 4587 19146 4597
rect 19272 4587 19338 4597
rect 19464 4587 19530 4597
rect 19656 4587 19722 4597
rect 20140 4587 20206 4597
rect 20332 4587 20398 4597
rect 20524 4587 20590 4597
rect 20716 4587 20782 4597
rect 20908 4587 20974 4597
rect 21100 4587 21166 4597
rect 21292 4587 21358 4597
rect 21484 4587 21550 4597
rect 128 4537 194 4547
rect 320 4537 386 4547
rect 512 4537 578 4547
rect 704 4537 770 4547
rect 896 4537 962 4547
rect 1088 4537 1154 4547
rect 1280 4537 1346 4547
rect 1472 4537 1528 4547
rect 1956 4537 2022 4547
rect 2148 4537 2214 4547
rect 2340 4537 2406 4547
rect 2532 4537 2598 4547
rect 2724 4537 2790 4547
rect 2916 4537 2982 4547
rect 3108 4537 3174 4547
rect 3300 4537 3356 4547
rect 3784 4537 3850 4547
rect 3976 4537 4042 4547
rect 4168 4537 4234 4547
rect 4360 4537 4426 4547
rect 4552 4537 4618 4547
rect 4744 4537 4810 4547
rect 4936 4537 5002 4547
rect 5128 4537 5184 4547
rect 5612 4537 5678 4547
rect 5804 4537 5870 4547
rect 5996 4537 6062 4547
rect 6188 4537 6254 4547
rect 6380 4537 6446 4547
rect 6572 4537 6638 4547
rect 6764 4537 6830 4547
rect 6956 4537 7012 4547
rect 7440 4537 7506 4547
rect 7632 4537 7698 4547
rect 7824 4537 7890 4547
rect 8016 4537 8082 4547
rect 8208 4537 8274 4547
rect 8400 4537 8466 4547
rect 8592 4537 8658 4547
rect 8784 4537 8840 4547
rect 9268 4537 9334 4547
rect 9460 4537 9526 4547
rect 9652 4537 9718 4547
rect 9844 4537 9910 4547
rect 10036 4537 10102 4547
rect 10228 4537 10294 4547
rect 10420 4537 10486 4547
rect 10612 4537 10668 4547
rect 11096 4537 11162 4547
rect 11288 4537 11354 4547
rect 11480 4537 11546 4547
rect 11672 4537 11738 4547
rect 11864 4537 11930 4547
rect 12056 4537 12122 4547
rect 12248 4537 12314 4547
rect 12440 4537 12496 4547
rect 12924 4537 12990 4547
rect 13116 4537 13182 4547
rect 13308 4537 13374 4547
rect 13500 4537 13566 4547
rect 13692 4537 13758 4547
rect 13884 4537 13950 4547
rect 14076 4537 14142 4547
rect 14268 4537 14324 4547
rect 14752 4537 14818 4547
rect 14944 4537 15010 4547
rect 15136 4537 15202 4547
rect 15328 4537 15394 4547
rect 15520 4537 15586 4547
rect 15712 4537 15778 4547
rect 15904 4537 15970 4547
rect 16096 4537 16152 4547
rect 16580 4537 16646 4547
rect 16772 4537 16838 4547
rect 16964 4537 17030 4547
rect 17156 4537 17222 4547
rect 17348 4537 17414 4547
rect 17540 4537 17606 4547
rect 17732 4537 17798 4547
rect 17924 4537 17980 4547
rect 18408 4537 18474 4547
rect 18600 4537 18666 4547
rect 18792 4537 18858 4547
rect 18984 4537 19050 4547
rect 19176 4537 19242 4547
rect 19368 4537 19434 4547
rect 19560 4537 19626 4547
rect 19752 4537 19808 4547
rect 20236 4537 20302 4547
rect 20428 4537 20494 4547
rect 20620 4537 20686 4547
rect 20812 4537 20878 4547
rect 21004 4537 21070 4547
rect 21196 4537 21262 4547
rect 21388 4537 21454 4547
rect 21580 4537 21636 4547
rect 0 4384 128 4537
rect 194 4384 320 4537
rect 386 4384 512 4537
rect 578 4384 704 4537
rect 770 4384 896 4537
rect 962 4384 1088 4537
rect 1154 4384 1280 4537
rect 1346 4384 1472 4537
rect 1528 4384 1708 4537
rect 1828 4384 1956 4537
rect 2022 4384 2148 4537
rect 2214 4384 2340 4537
rect 2406 4384 2532 4537
rect 2598 4384 2724 4537
rect 2790 4384 2916 4537
rect 2982 4384 3108 4537
rect 3174 4384 3300 4537
rect 3356 4384 3536 4537
rect 3656 4384 3784 4537
rect 3850 4384 3976 4537
rect 4042 4384 4168 4537
rect 4234 4384 4360 4537
rect 4426 4384 4552 4537
rect 4618 4384 4744 4537
rect 4810 4384 4936 4537
rect 5002 4384 5128 4537
rect 5184 4384 5364 4537
rect 5484 4384 5612 4537
rect 5678 4384 5804 4537
rect 5870 4384 5996 4537
rect 6062 4384 6188 4537
rect 6254 4384 6380 4537
rect 6446 4384 6572 4537
rect 6638 4384 6764 4537
rect 6830 4384 6956 4537
rect 7012 4384 7192 4537
rect 7312 4384 7440 4537
rect 7506 4384 7632 4537
rect 7698 4384 7824 4537
rect 7890 4384 8016 4537
rect 8082 4384 8208 4537
rect 8274 4384 8400 4537
rect 8466 4384 8592 4537
rect 8658 4384 8784 4537
rect 8840 4384 9020 4537
rect 9140 4384 9268 4537
rect 9334 4384 9460 4537
rect 9526 4384 9652 4537
rect 9718 4384 9844 4537
rect 9910 4384 10036 4537
rect 10102 4384 10228 4537
rect 10294 4384 10420 4537
rect 10486 4384 10612 4537
rect 10668 4384 10848 4537
rect 10968 4384 11096 4537
rect 11162 4384 11288 4537
rect 11354 4384 11480 4537
rect 11546 4384 11672 4537
rect 11738 4384 11864 4537
rect 11930 4384 12056 4537
rect 12122 4384 12248 4537
rect 12314 4384 12440 4537
rect 12496 4384 12676 4537
rect 12796 4384 12924 4537
rect 12990 4384 13116 4537
rect 13182 4384 13308 4537
rect 13374 4384 13500 4537
rect 13566 4384 13692 4537
rect 13758 4384 13884 4537
rect 13950 4384 14076 4537
rect 14142 4384 14268 4537
rect 14324 4384 14504 4537
rect 14624 4384 14752 4537
rect 14818 4384 14944 4537
rect 15010 4384 15136 4537
rect 15202 4384 15328 4537
rect 15394 4384 15520 4537
rect 15586 4384 15712 4537
rect 15778 4384 15904 4537
rect 15970 4384 16096 4537
rect 16152 4384 16332 4537
rect 16452 4384 16580 4537
rect 16646 4384 16772 4537
rect 16838 4384 16964 4537
rect 17030 4384 17156 4537
rect 17222 4384 17348 4537
rect 17414 4384 17540 4537
rect 17606 4384 17732 4537
rect 17798 4384 17924 4537
rect 17980 4384 18160 4537
rect 18280 4384 18408 4537
rect 18474 4384 18600 4537
rect 18666 4384 18792 4537
rect 18858 4384 18984 4537
rect 19050 4384 19176 4537
rect 19242 4384 19368 4537
rect 19434 4384 19560 4537
rect 19626 4384 19752 4537
rect 19808 4384 19988 4537
rect 20108 4384 20236 4537
rect 20302 4384 20428 4537
rect 20494 4384 20620 4537
rect 20686 4384 20812 4537
rect 20878 4384 21004 4537
rect 21070 4384 21196 4537
rect 21262 4384 21388 4537
rect 21454 4384 21580 4537
rect 21636 4384 21816 4537
rect 128 4374 194 4384
rect 320 4374 386 4384
rect 512 4374 578 4384
rect 704 4374 770 4384
rect 896 4374 962 4384
rect 1088 4374 1154 4384
rect 1280 4374 1346 4384
rect 1472 4374 1528 4384
rect 1956 4374 2022 4384
rect 2148 4374 2214 4384
rect 2340 4374 2406 4384
rect 2532 4374 2598 4384
rect 2724 4374 2790 4384
rect 2916 4374 2982 4384
rect 3108 4374 3174 4384
rect 3300 4374 3356 4384
rect 3784 4374 3850 4384
rect 3976 4374 4042 4384
rect 4168 4374 4234 4384
rect 4360 4374 4426 4384
rect 4552 4374 4618 4384
rect 4744 4374 4810 4384
rect 4936 4374 5002 4384
rect 5128 4374 5184 4384
rect 5612 4374 5678 4384
rect 5804 4374 5870 4384
rect 5996 4374 6062 4384
rect 6188 4374 6254 4384
rect 6380 4374 6446 4384
rect 6572 4374 6638 4384
rect 6764 4374 6830 4384
rect 6956 4374 7012 4384
rect 7440 4374 7506 4384
rect 7632 4374 7698 4384
rect 7824 4374 7890 4384
rect 8016 4374 8082 4384
rect 8208 4374 8274 4384
rect 8400 4374 8466 4384
rect 8592 4374 8658 4384
rect 8784 4374 8840 4384
rect 9268 4374 9334 4384
rect 9460 4374 9526 4384
rect 9652 4374 9718 4384
rect 9844 4374 9910 4384
rect 10036 4374 10102 4384
rect 10228 4374 10294 4384
rect 10420 4374 10486 4384
rect 10612 4374 10668 4384
rect 11096 4374 11162 4384
rect 11288 4374 11354 4384
rect 11480 4374 11546 4384
rect 11672 4374 11738 4384
rect 11864 4374 11930 4384
rect 12056 4374 12122 4384
rect 12248 4374 12314 4384
rect 12440 4374 12496 4384
rect 12924 4374 12990 4384
rect 13116 4374 13182 4384
rect 13308 4374 13374 4384
rect 13500 4374 13566 4384
rect 13692 4374 13758 4384
rect 13884 4374 13950 4384
rect 14076 4374 14142 4384
rect 14268 4374 14324 4384
rect 14752 4374 14818 4384
rect 14944 4374 15010 4384
rect 15136 4374 15202 4384
rect 15328 4374 15394 4384
rect 15520 4374 15586 4384
rect 15712 4374 15778 4384
rect 15904 4374 15970 4384
rect 16096 4374 16152 4384
rect 16580 4374 16646 4384
rect 16772 4374 16838 4384
rect 16964 4374 17030 4384
rect 17156 4374 17222 4384
rect 17348 4374 17414 4384
rect 17540 4374 17606 4384
rect 17732 4374 17798 4384
rect 17924 4374 17980 4384
rect 18408 4374 18474 4384
rect 18600 4374 18666 4384
rect 18792 4374 18858 4384
rect 18984 4374 19050 4384
rect 19176 4374 19242 4384
rect 19368 4374 19434 4384
rect 19560 4374 19626 4384
rect 19752 4374 19808 4384
rect 20236 4374 20302 4384
rect 20428 4374 20494 4384
rect 20620 4374 20686 4384
rect 20812 4374 20878 4384
rect 21004 4374 21070 4384
rect 21196 4374 21262 4384
rect 21388 4374 21454 4384
rect 21580 4374 21636 4384
rect 32 4036 98 4046
rect 224 4036 290 4046
rect 416 4036 482 4046
rect 608 4036 674 4046
rect 800 4036 866 4046
rect 992 4036 1058 4046
rect 1184 4036 1250 4046
rect 1376 4036 1442 4046
rect 1860 4036 1926 4046
rect 2052 4036 2118 4046
rect 2244 4036 2310 4046
rect 2436 4036 2502 4046
rect 2628 4036 2694 4046
rect 2820 4036 2886 4046
rect 3012 4036 3078 4046
rect 3204 4036 3270 4046
rect 3688 4036 3754 4046
rect 3880 4036 3946 4046
rect 4072 4036 4138 4046
rect 4264 4036 4330 4046
rect 4456 4036 4522 4046
rect 4648 4036 4714 4046
rect 4840 4036 4906 4046
rect 5032 4036 5098 4046
rect 5516 4036 5582 4046
rect 5708 4036 5774 4046
rect 5900 4036 5966 4046
rect 6092 4036 6158 4046
rect 6284 4036 6350 4046
rect 6476 4036 6542 4046
rect 6668 4036 6734 4046
rect 6860 4036 6926 4046
rect 7344 4036 7410 4046
rect 7536 4036 7602 4046
rect 7728 4036 7794 4046
rect 7920 4036 7986 4046
rect 8112 4036 8178 4046
rect 8304 4036 8370 4046
rect 8496 4036 8562 4046
rect 8688 4036 8754 4046
rect 9172 4036 9238 4046
rect 9364 4036 9430 4046
rect 9556 4036 9622 4046
rect 9748 4036 9814 4046
rect 9940 4036 10006 4046
rect 10132 4036 10198 4046
rect 10324 4036 10390 4046
rect 10516 4036 10582 4046
rect 11000 4036 11066 4046
rect 11192 4036 11258 4046
rect 11384 4036 11450 4046
rect 11576 4036 11642 4046
rect 11768 4036 11834 4046
rect 11960 4036 12026 4046
rect 12152 4036 12218 4046
rect 12344 4036 12410 4046
rect 12828 4036 12894 4046
rect 13020 4036 13086 4046
rect 13212 4036 13278 4046
rect 13404 4036 13470 4046
rect 13596 4036 13662 4046
rect 13788 4036 13854 4046
rect 13980 4036 14046 4046
rect 14172 4036 14238 4046
rect 14656 4036 14722 4046
rect 14848 4036 14914 4046
rect 15040 4036 15106 4046
rect 15232 4036 15298 4046
rect 15424 4036 15490 4046
rect 15616 4036 15682 4046
rect 15808 4036 15874 4046
rect 16000 4036 16066 4046
rect 16484 4036 16550 4046
rect 16676 4036 16742 4046
rect 16868 4036 16934 4046
rect 17060 4036 17126 4046
rect 17252 4036 17318 4046
rect 17444 4036 17510 4046
rect 17636 4036 17702 4046
rect 17828 4036 17894 4046
rect 18312 4036 18378 4046
rect 18504 4036 18570 4046
rect 18696 4036 18762 4046
rect 18888 4036 18954 4046
rect 19080 4036 19146 4046
rect 19272 4036 19338 4046
rect 19464 4036 19530 4046
rect 19656 4036 19722 4046
rect 20140 4036 20206 4046
rect 20332 4036 20398 4046
rect 20524 4036 20590 4046
rect 20716 4036 20782 4046
rect 20908 4036 20974 4046
rect 21100 4036 21166 4046
rect 21292 4036 21358 4046
rect 21484 4036 21550 4046
rect 0 3883 32 4036
rect 98 3883 224 4036
rect 290 3883 416 4036
rect 482 3883 608 4036
rect 674 3883 800 4036
rect 866 3883 992 4036
rect 1058 3883 1184 4036
rect 1250 3883 1376 4036
rect 1828 3883 1860 4036
rect 1926 3883 2052 4036
rect 2118 3883 2244 4036
rect 2310 3883 2436 4036
rect 2502 3883 2628 4036
rect 2694 3883 2820 4036
rect 2886 3883 3012 4036
rect 3078 3883 3204 4036
rect 3656 3883 3688 4036
rect 3754 3883 3880 4036
rect 3946 3883 4072 4036
rect 4138 3883 4264 4036
rect 4330 3883 4456 4036
rect 4522 3883 4648 4036
rect 4714 3883 4840 4036
rect 4906 3883 5032 4036
rect 5484 3883 5516 4036
rect 5582 3883 5708 4036
rect 5774 3883 5900 4036
rect 5966 3883 6092 4036
rect 6158 3883 6284 4036
rect 6350 3883 6476 4036
rect 6542 3883 6668 4036
rect 6734 3883 6860 4036
rect 7312 3883 7344 4036
rect 7410 3883 7536 4036
rect 7602 3883 7728 4036
rect 7794 3883 7920 4036
rect 7986 3883 8112 4036
rect 8178 3883 8304 4036
rect 8370 3883 8496 4036
rect 8562 3883 8688 4036
rect 9140 3883 9172 4036
rect 9238 3883 9364 4036
rect 9430 3883 9556 4036
rect 9622 3883 9748 4036
rect 9814 3883 9940 4036
rect 10006 3883 10132 4036
rect 10198 3883 10324 4036
rect 10390 3883 10516 4036
rect 10968 3883 11000 4036
rect 11066 3883 11192 4036
rect 11258 3883 11384 4036
rect 11450 3883 11576 4036
rect 11642 3883 11768 4036
rect 11834 3883 11960 4036
rect 12026 3883 12152 4036
rect 12218 3883 12344 4036
rect 12796 3883 12828 4036
rect 12894 3883 13020 4036
rect 13086 3883 13212 4036
rect 13278 3883 13404 4036
rect 13470 3883 13596 4036
rect 13662 3883 13788 4036
rect 13854 3883 13980 4036
rect 14046 3883 14172 4036
rect 14624 3883 14656 4036
rect 14722 3883 14848 4036
rect 14914 3883 15040 4036
rect 15106 3883 15232 4036
rect 15298 3883 15424 4036
rect 15490 3883 15616 4036
rect 15682 3883 15808 4036
rect 15874 3883 16000 4036
rect 16452 3883 16484 4036
rect 16550 3883 16676 4036
rect 16742 3883 16868 4036
rect 16934 3883 17060 4036
rect 17126 3883 17252 4036
rect 17318 3883 17444 4036
rect 17510 3883 17636 4036
rect 17702 3883 17828 4036
rect 18280 3883 18312 4036
rect 18378 3883 18504 4036
rect 18570 3883 18696 4036
rect 18762 3883 18888 4036
rect 18954 3883 19080 4036
rect 19146 3883 19272 4036
rect 19338 3883 19464 4036
rect 19530 3883 19656 4036
rect 20108 3883 20140 4036
rect 20206 3883 20332 4036
rect 20398 3883 20524 4036
rect 20590 3883 20716 4036
rect 20782 3883 20908 4036
rect 20974 3883 21100 4036
rect 21166 3883 21292 4036
rect 21358 3883 21484 4036
rect 32 3873 98 3883
rect 224 3873 290 3883
rect 416 3873 482 3883
rect 608 3873 674 3883
rect 800 3873 866 3883
rect 992 3873 1058 3883
rect 1184 3873 1250 3883
rect 1376 3873 1442 3883
rect 1860 3873 1926 3883
rect 2052 3873 2118 3883
rect 2244 3873 2310 3883
rect 2436 3873 2502 3883
rect 2628 3873 2694 3883
rect 2820 3873 2886 3883
rect 3012 3873 3078 3883
rect 3204 3873 3270 3883
rect 3688 3873 3754 3883
rect 3880 3873 3946 3883
rect 4072 3873 4138 3883
rect 4264 3873 4330 3883
rect 4456 3873 4522 3883
rect 4648 3873 4714 3883
rect 4840 3873 4906 3883
rect 5032 3873 5098 3883
rect 5516 3873 5582 3883
rect 5708 3873 5774 3883
rect 5900 3873 5966 3883
rect 6092 3873 6158 3883
rect 6284 3873 6350 3883
rect 6476 3873 6542 3883
rect 6668 3873 6734 3883
rect 6860 3873 6926 3883
rect 7344 3873 7410 3883
rect 7536 3873 7602 3883
rect 7728 3873 7794 3883
rect 7920 3873 7986 3883
rect 8112 3873 8178 3883
rect 8304 3873 8370 3883
rect 8496 3873 8562 3883
rect 8688 3873 8754 3883
rect 9172 3873 9238 3883
rect 9364 3873 9430 3883
rect 9556 3873 9622 3883
rect 9748 3873 9814 3883
rect 9940 3873 10006 3883
rect 10132 3873 10198 3883
rect 10324 3873 10390 3883
rect 10516 3873 10582 3883
rect 11000 3873 11066 3883
rect 11192 3873 11258 3883
rect 11384 3873 11450 3883
rect 11576 3873 11642 3883
rect 11768 3873 11834 3883
rect 11960 3873 12026 3883
rect 12152 3873 12218 3883
rect 12344 3873 12410 3883
rect 12828 3873 12894 3883
rect 13020 3873 13086 3883
rect 13212 3873 13278 3883
rect 13404 3873 13470 3883
rect 13596 3873 13662 3883
rect 13788 3873 13854 3883
rect 13980 3873 14046 3883
rect 14172 3873 14238 3883
rect 14656 3873 14722 3883
rect 14848 3873 14914 3883
rect 15040 3873 15106 3883
rect 15232 3873 15298 3883
rect 15424 3873 15490 3883
rect 15616 3873 15682 3883
rect 15808 3873 15874 3883
rect 16000 3873 16066 3883
rect 16484 3873 16550 3883
rect 16676 3873 16742 3883
rect 16868 3873 16934 3883
rect 17060 3873 17126 3883
rect 17252 3873 17318 3883
rect 17444 3873 17510 3883
rect 17636 3873 17702 3883
rect 17828 3873 17894 3883
rect 18312 3873 18378 3883
rect 18504 3873 18570 3883
rect 18696 3873 18762 3883
rect 18888 3873 18954 3883
rect 19080 3873 19146 3883
rect 19272 3873 19338 3883
rect 19464 3873 19530 3883
rect 19656 3873 19722 3883
rect 20140 3873 20206 3883
rect 20332 3873 20398 3883
rect 20524 3873 20590 3883
rect 20716 3873 20782 3883
rect 20908 3873 20974 3883
rect 21100 3873 21166 3883
rect 21292 3873 21358 3883
rect 21484 3873 21550 3883
rect 128 3823 194 3833
rect 320 3823 386 3833
rect 512 3823 578 3833
rect 704 3823 770 3833
rect 896 3823 962 3833
rect 1088 3823 1154 3833
rect 1280 3823 1346 3833
rect 1472 3823 1528 3833
rect 1956 3823 2022 3833
rect 2148 3823 2214 3833
rect 2340 3823 2406 3833
rect 2532 3823 2598 3833
rect 2724 3823 2790 3833
rect 2916 3823 2982 3833
rect 3108 3823 3174 3833
rect 3300 3823 3356 3833
rect 3784 3823 3850 3833
rect 3976 3823 4042 3833
rect 4168 3823 4234 3833
rect 4360 3823 4426 3833
rect 4552 3823 4618 3833
rect 4744 3823 4810 3833
rect 4936 3823 5002 3833
rect 5128 3823 5184 3833
rect 5612 3823 5678 3833
rect 5804 3823 5870 3833
rect 5996 3823 6062 3833
rect 6188 3823 6254 3833
rect 6380 3823 6446 3833
rect 6572 3823 6638 3833
rect 6764 3823 6830 3833
rect 6956 3823 7012 3833
rect 7440 3823 7506 3833
rect 7632 3823 7698 3833
rect 7824 3823 7890 3833
rect 8016 3823 8082 3833
rect 8208 3823 8274 3833
rect 8400 3823 8466 3833
rect 8592 3823 8658 3833
rect 8784 3823 8840 3833
rect 9268 3823 9334 3833
rect 9460 3823 9526 3833
rect 9652 3823 9718 3833
rect 9844 3823 9910 3833
rect 10036 3823 10102 3833
rect 10228 3823 10294 3833
rect 10420 3823 10486 3833
rect 10612 3823 10668 3833
rect 11096 3823 11162 3833
rect 11288 3823 11354 3833
rect 11480 3823 11546 3833
rect 11672 3823 11738 3833
rect 11864 3823 11930 3833
rect 12056 3823 12122 3833
rect 12248 3823 12314 3833
rect 12440 3823 12496 3833
rect 12924 3823 12990 3833
rect 13116 3823 13182 3833
rect 13308 3823 13374 3833
rect 13500 3823 13566 3833
rect 13692 3823 13758 3833
rect 13884 3823 13950 3833
rect 14076 3823 14142 3833
rect 14268 3823 14324 3833
rect 14752 3823 14818 3833
rect 14944 3823 15010 3833
rect 15136 3823 15202 3833
rect 15328 3823 15394 3833
rect 15520 3823 15586 3833
rect 15712 3823 15778 3833
rect 15904 3823 15970 3833
rect 16096 3823 16152 3833
rect 16580 3823 16646 3833
rect 16772 3823 16838 3833
rect 16964 3823 17030 3833
rect 17156 3823 17222 3833
rect 17348 3823 17414 3833
rect 17540 3823 17606 3833
rect 17732 3823 17798 3833
rect 17924 3823 17980 3833
rect 18408 3823 18474 3833
rect 18600 3823 18666 3833
rect 18792 3823 18858 3833
rect 18984 3823 19050 3833
rect 19176 3823 19242 3833
rect 19368 3823 19434 3833
rect 19560 3823 19626 3833
rect 19752 3823 19808 3833
rect 20236 3823 20302 3833
rect 20428 3823 20494 3833
rect 20620 3823 20686 3833
rect 20812 3823 20878 3833
rect 21004 3823 21070 3833
rect 21196 3823 21262 3833
rect 21388 3823 21454 3833
rect 21580 3823 21636 3833
rect 0 3670 128 3823
rect 194 3670 320 3823
rect 386 3670 512 3823
rect 578 3670 704 3823
rect 770 3670 896 3823
rect 962 3670 1088 3823
rect 1154 3670 1280 3823
rect 1346 3670 1472 3823
rect 1528 3670 1708 3823
rect 1828 3670 1956 3823
rect 2022 3670 2148 3823
rect 2214 3670 2340 3823
rect 2406 3670 2532 3823
rect 2598 3670 2724 3823
rect 2790 3670 2916 3823
rect 2982 3670 3108 3823
rect 3174 3670 3300 3823
rect 3356 3670 3536 3823
rect 3656 3670 3784 3823
rect 3850 3670 3976 3823
rect 4042 3670 4168 3823
rect 4234 3670 4360 3823
rect 4426 3670 4552 3823
rect 4618 3670 4744 3823
rect 4810 3670 4936 3823
rect 5002 3670 5128 3823
rect 5184 3670 5364 3823
rect 5484 3670 5612 3823
rect 5678 3670 5804 3823
rect 5870 3670 5996 3823
rect 6062 3670 6188 3823
rect 6254 3670 6380 3823
rect 6446 3670 6572 3823
rect 6638 3670 6764 3823
rect 6830 3670 6956 3823
rect 7012 3670 7192 3823
rect 7312 3670 7440 3823
rect 7506 3670 7632 3823
rect 7698 3670 7824 3823
rect 7890 3670 8016 3823
rect 8082 3670 8208 3823
rect 8274 3670 8400 3823
rect 8466 3670 8592 3823
rect 8658 3670 8784 3823
rect 8840 3670 9020 3823
rect 9140 3670 9268 3823
rect 9334 3670 9460 3823
rect 9526 3670 9652 3823
rect 9718 3670 9844 3823
rect 9910 3670 10036 3823
rect 10102 3670 10228 3823
rect 10294 3670 10420 3823
rect 10486 3670 10612 3823
rect 10668 3670 10848 3823
rect 10968 3670 11096 3823
rect 11162 3670 11288 3823
rect 11354 3670 11480 3823
rect 11546 3670 11672 3823
rect 11738 3670 11864 3823
rect 11930 3670 12056 3823
rect 12122 3670 12248 3823
rect 12314 3670 12440 3823
rect 12496 3670 12676 3823
rect 12796 3670 12924 3823
rect 12990 3670 13116 3823
rect 13182 3670 13308 3823
rect 13374 3670 13500 3823
rect 13566 3670 13692 3823
rect 13758 3670 13884 3823
rect 13950 3670 14076 3823
rect 14142 3670 14268 3823
rect 14324 3670 14504 3823
rect 14624 3670 14752 3823
rect 14818 3670 14944 3823
rect 15010 3670 15136 3823
rect 15202 3670 15328 3823
rect 15394 3670 15520 3823
rect 15586 3670 15712 3823
rect 15778 3670 15904 3823
rect 15970 3670 16096 3823
rect 16152 3670 16332 3823
rect 16452 3670 16580 3823
rect 16646 3670 16772 3823
rect 16838 3670 16964 3823
rect 17030 3670 17156 3823
rect 17222 3670 17348 3823
rect 17414 3670 17540 3823
rect 17606 3670 17732 3823
rect 17798 3670 17924 3823
rect 17980 3670 18160 3823
rect 18280 3670 18408 3823
rect 18474 3670 18600 3823
rect 18666 3670 18792 3823
rect 18858 3670 18984 3823
rect 19050 3670 19176 3823
rect 19242 3670 19368 3823
rect 19434 3670 19560 3823
rect 19626 3670 19752 3823
rect 19808 3670 19988 3823
rect 20108 3670 20236 3823
rect 20302 3670 20428 3823
rect 20494 3670 20620 3823
rect 20686 3670 20812 3823
rect 20878 3670 21004 3823
rect 21070 3670 21196 3823
rect 21262 3670 21388 3823
rect 21454 3670 21580 3823
rect 21636 3670 21816 3823
rect 128 3660 194 3670
rect 320 3660 386 3670
rect 512 3660 578 3670
rect 704 3660 770 3670
rect 896 3660 962 3670
rect 1088 3660 1154 3670
rect 1280 3660 1346 3670
rect 1472 3660 1528 3670
rect 1956 3660 2022 3670
rect 2148 3660 2214 3670
rect 2340 3660 2406 3670
rect 2532 3660 2598 3670
rect 2724 3660 2790 3670
rect 2916 3660 2982 3670
rect 3108 3660 3174 3670
rect 3300 3660 3356 3670
rect 3784 3660 3850 3670
rect 3976 3660 4042 3670
rect 4168 3660 4234 3670
rect 4360 3660 4426 3670
rect 4552 3660 4618 3670
rect 4744 3660 4810 3670
rect 4936 3660 5002 3670
rect 5128 3660 5184 3670
rect 5612 3660 5678 3670
rect 5804 3660 5870 3670
rect 5996 3660 6062 3670
rect 6188 3660 6254 3670
rect 6380 3660 6446 3670
rect 6572 3660 6638 3670
rect 6764 3660 6830 3670
rect 6956 3660 7012 3670
rect 7440 3660 7506 3670
rect 7632 3660 7698 3670
rect 7824 3660 7890 3670
rect 8016 3660 8082 3670
rect 8208 3660 8274 3670
rect 8400 3660 8466 3670
rect 8592 3660 8658 3670
rect 8784 3660 8840 3670
rect 9268 3660 9334 3670
rect 9460 3660 9526 3670
rect 9652 3660 9718 3670
rect 9844 3660 9910 3670
rect 10036 3660 10102 3670
rect 10228 3660 10294 3670
rect 10420 3660 10486 3670
rect 10612 3660 10668 3670
rect 11096 3660 11162 3670
rect 11288 3660 11354 3670
rect 11480 3660 11546 3670
rect 11672 3660 11738 3670
rect 11864 3660 11930 3670
rect 12056 3660 12122 3670
rect 12248 3660 12314 3670
rect 12440 3660 12496 3670
rect 12924 3660 12990 3670
rect 13116 3660 13182 3670
rect 13308 3660 13374 3670
rect 13500 3660 13566 3670
rect 13692 3660 13758 3670
rect 13884 3660 13950 3670
rect 14076 3660 14142 3670
rect 14268 3660 14324 3670
rect 14752 3660 14818 3670
rect 14944 3660 15010 3670
rect 15136 3660 15202 3670
rect 15328 3660 15394 3670
rect 15520 3660 15586 3670
rect 15712 3660 15778 3670
rect 15904 3660 15970 3670
rect 16096 3660 16152 3670
rect 16580 3660 16646 3670
rect 16772 3660 16838 3670
rect 16964 3660 17030 3670
rect 17156 3660 17222 3670
rect 17348 3660 17414 3670
rect 17540 3660 17606 3670
rect 17732 3660 17798 3670
rect 17924 3660 17980 3670
rect 18408 3660 18474 3670
rect 18600 3660 18666 3670
rect 18792 3660 18858 3670
rect 18984 3660 19050 3670
rect 19176 3660 19242 3670
rect 19368 3660 19434 3670
rect 19560 3660 19626 3670
rect 19752 3660 19808 3670
rect 20236 3660 20302 3670
rect 20428 3660 20494 3670
rect 20620 3660 20686 3670
rect 20812 3660 20878 3670
rect 21004 3660 21070 3670
rect 21196 3660 21262 3670
rect 21388 3660 21454 3670
rect 21580 3660 21636 3670
rect 32 3322 98 3332
rect 224 3322 290 3332
rect 416 3322 482 3332
rect 608 3322 674 3332
rect 800 3322 866 3332
rect 992 3322 1058 3332
rect 1184 3322 1250 3332
rect 1376 3322 1442 3332
rect 1860 3322 1926 3332
rect 2052 3322 2118 3332
rect 2244 3322 2310 3332
rect 2436 3322 2502 3332
rect 2628 3322 2694 3332
rect 2820 3322 2886 3332
rect 3012 3322 3078 3332
rect 3204 3322 3270 3332
rect 3688 3322 3754 3332
rect 3880 3322 3946 3332
rect 4072 3322 4138 3332
rect 4264 3322 4330 3332
rect 4456 3322 4522 3332
rect 4648 3322 4714 3332
rect 4840 3322 4906 3332
rect 5032 3322 5098 3332
rect 5516 3322 5582 3332
rect 5708 3322 5774 3332
rect 5900 3322 5966 3332
rect 6092 3322 6158 3332
rect 6284 3322 6350 3332
rect 6476 3322 6542 3332
rect 6668 3322 6734 3332
rect 6860 3322 6926 3332
rect 7344 3322 7410 3332
rect 7536 3322 7602 3332
rect 7728 3322 7794 3332
rect 7920 3322 7986 3332
rect 8112 3322 8178 3332
rect 8304 3322 8370 3332
rect 8496 3322 8562 3332
rect 8688 3322 8754 3332
rect 9172 3322 9238 3332
rect 9364 3322 9430 3332
rect 9556 3322 9622 3332
rect 9748 3322 9814 3332
rect 9940 3322 10006 3332
rect 10132 3322 10198 3332
rect 10324 3322 10390 3332
rect 10516 3322 10582 3332
rect 11000 3322 11066 3332
rect 11192 3322 11258 3332
rect 11384 3322 11450 3332
rect 11576 3322 11642 3332
rect 11768 3322 11834 3332
rect 11960 3322 12026 3332
rect 12152 3322 12218 3332
rect 12344 3322 12410 3332
rect 12828 3322 12894 3332
rect 13020 3322 13086 3332
rect 13212 3322 13278 3332
rect 13404 3322 13470 3332
rect 13596 3322 13662 3332
rect 13788 3322 13854 3332
rect 13980 3322 14046 3332
rect 14172 3322 14238 3332
rect 14656 3322 14722 3332
rect 14848 3322 14914 3332
rect 15040 3322 15106 3332
rect 15232 3322 15298 3332
rect 15424 3322 15490 3332
rect 15616 3322 15682 3332
rect 15808 3322 15874 3332
rect 16000 3322 16066 3332
rect 16484 3322 16550 3332
rect 16676 3322 16742 3332
rect 16868 3322 16934 3332
rect 17060 3322 17126 3332
rect 17252 3322 17318 3332
rect 17444 3322 17510 3332
rect 17636 3322 17702 3332
rect 17828 3322 17894 3332
rect 18312 3322 18378 3332
rect 18504 3322 18570 3332
rect 18696 3322 18762 3332
rect 18888 3322 18954 3332
rect 19080 3322 19146 3332
rect 19272 3322 19338 3332
rect 19464 3322 19530 3332
rect 19656 3322 19722 3332
rect 20140 3322 20206 3332
rect 20332 3322 20398 3332
rect 20524 3322 20590 3332
rect 20716 3322 20782 3332
rect 20908 3322 20974 3332
rect 21100 3322 21166 3332
rect 21292 3322 21358 3332
rect 21484 3322 21550 3332
rect 0 3169 32 3322
rect 98 3169 224 3322
rect 290 3169 416 3322
rect 482 3169 608 3322
rect 674 3169 800 3322
rect 866 3169 992 3322
rect 1058 3169 1184 3322
rect 1250 3169 1376 3322
rect 1828 3169 1860 3322
rect 1926 3169 2052 3322
rect 2118 3169 2244 3322
rect 2310 3169 2436 3322
rect 2502 3169 2628 3322
rect 2694 3169 2820 3322
rect 2886 3169 3012 3322
rect 3078 3169 3204 3322
rect 3656 3169 3688 3322
rect 3754 3169 3880 3322
rect 3946 3169 4072 3322
rect 4138 3169 4264 3322
rect 4330 3169 4456 3322
rect 4522 3169 4648 3322
rect 4714 3169 4840 3322
rect 4906 3169 5032 3322
rect 5484 3169 5516 3322
rect 5582 3169 5708 3322
rect 5774 3169 5900 3322
rect 5966 3169 6092 3322
rect 6158 3169 6284 3322
rect 6350 3169 6476 3322
rect 6542 3169 6668 3322
rect 6734 3169 6860 3322
rect 7312 3169 7344 3322
rect 7410 3169 7536 3322
rect 7602 3169 7728 3322
rect 7794 3169 7920 3322
rect 7986 3169 8112 3322
rect 8178 3169 8304 3322
rect 8370 3169 8496 3322
rect 8562 3169 8688 3322
rect 9140 3169 9172 3322
rect 9238 3169 9364 3322
rect 9430 3169 9556 3322
rect 9622 3169 9748 3322
rect 9814 3169 9940 3322
rect 10006 3169 10132 3322
rect 10198 3169 10324 3322
rect 10390 3169 10516 3322
rect 10968 3169 11000 3322
rect 11066 3169 11192 3322
rect 11258 3169 11384 3322
rect 11450 3169 11576 3322
rect 11642 3169 11768 3322
rect 11834 3169 11960 3322
rect 12026 3169 12152 3322
rect 12218 3169 12344 3322
rect 12796 3169 12828 3322
rect 12894 3169 13020 3322
rect 13086 3169 13212 3322
rect 13278 3169 13404 3322
rect 13470 3169 13596 3322
rect 13662 3169 13788 3322
rect 13854 3169 13980 3322
rect 14046 3169 14172 3322
rect 14624 3169 14656 3322
rect 14722 3169 14848 3322
rect 14914 3169 15040 3322
rect 15106 3169 15232 3322
rect 15298 3169 15424 3322
rect 15490 3169 15616 3322
rect 15682 3169 15808 3322
rect 15874 3169 16000 3322
rect 16452 3169 16484 3322
rect 16550 3169 16676 3322
rect 16742 3169 16868 3322
rect 16934 3169 17060 3322
rect 17126 3169 17252 3322
rect 17318 3169 17444 3322
rect 17510 3169 17636 3322
rect 17702 3169 17828 3322
rect 18280 3169 18312 3322
rect 18378 3169 18504 3322
rect 18570 3169 18696 3322
rect 18762 3169 18888 3322
rect 18954 3169 19080 3322
rect 19146 3169 19272 3322
rect 19338 3169 19464 3322
rect 19530 3169 19656 3322
rect 20108 3169 20140 3322
rect 20206 3169 20332 3322
rect 20398 3169 20524 3322
rect 20590 3169 20716 3322
rect 20782 3169 20908 3322
rect 20974 3169 21100 3322
rect 21166 3169 21292 3322
rect 21358 3169 21484 3322
rect 32 3159 98 3169
rect 224 3159 290 3169
rect 416 3159 482 3169
rect 608 3159 674 3169
rect 800 3159 866 3169
rect 992 3159 1058 3169
rect 1184 3159 1250 3169
rect 1376 3159 1442 3169
rect 1860 3159 1926 3169
rect 2052 3159 2118 3169
rect 2244 3159 2310 3169
rect 2436 3159 2502 3169
rect 2628 3159 2694 3169
rect 2820 3159 2886 3169
rect 3012 3159 3078 3169
rect 3204 3159 3270 3169
rect 3688 3159 3754 3169
rect 3880 3159 3946 3169
rect 4072 3159 4138 3169
rect 4264 3159 4330 3169
rect 4456 3159 4522 3169
rect 4648 3159 4714 3169
rect 4840 3159 4906 3169
rect 5032 3159 5098 3169
rect 5516 3159 5582 3169
rect 5708 3159 5774 3169
rect 5900 3159 5966 3169
rect 6092 3159 6158 3169
rect 6284 3159 6350 3169
rect 6476 3159 6542 3169
rect 6668 3159 6734 3169
rect 6860 3159 6926 3169
rect 7344 3159 7410 3169
rect 7536 3159 7602 3169
rect 7728 3159 7794 3169
rect 7920 3159 7986 3169
rect 8112 3159 8178 3169
rect 8304 3159 8370 3169
rect 8496 3159 8562 3169
rect 8688 3159 8754 3169
rect 9172 3159 9238 3169
rect 9364 3159 9430 3169
rect 9556 3159 9622 3169
rect 9748 3159 9814 3169
rect 9940 3159 10006 3169
rect 10132 3159 10198 3169
rect 10324 3159 10390 3169
rect 10516 3159 10582 3169
rect 11000 3159 11066 3169
rect 11192 3159 11258 3169
rect 11384 3159 11450 3169
rect 11576 3159 11642 3169
rect 11768 3159 11834 3169
rect 11960 3159 12026 3169
rect 12152 3159 12218 3169
rect 12344 3159 12410 3169
rect 12828 3159 12894 3169
rect 13020 3159 13086 3169
rect 13212 3159 13278 3169
rect 13404 3159 13470 3169
rect 13596 3159 13662 3169
rect 13788 3159 13854 3169
rect 13980 3159 14046 3169
rect 14172 3159 14238 3169
rect 14656 3159 14722 3169
rect 14848 3159 14914 3169
rect 15040 3159 15106 3169
rect 15232 3159 15298 3169
rect 15424 3159 15490 3169
rect 15616 3159 15682 3169
rect 15808 3159 15874 3169
rect 16000 3159 16066 3169
rect 16484 3159 16550 3169
rect 16676 3159 16742 3169
rect 16868 3159 16934 3169
rect 17060 3159 17126 3169
rect 17252 3159 17318 3169
rect 17444 3159 17510 3169
rect 17636 3159 17702 3169
rect 17828 3159 17894 3169
rect 18312 3159 18378 3169
rect 18504 3159 18570 3169
rect 18696 3159 18762 3169
rect 18888 3159 18954 3169
rect 19080 3159 19146 3169
rect 19272 3159 19338 3169
rect 19464 3159 19530 3169
rect 19656 3159 19722 3169
rect 20140 3159 20206 3169
rect 20332 3159 20398 3169
rect 20524 3159 20590 3169
rect 20716 3159 20782 3169
rect 20908 3159 20974 3169
rect 21100 3159 21166 3169
rect 21292 3159 21358 3169
rect 21484 3159 21550 3169
rect 128 3109 194 3119
rect 320 3109 386 3119
rect 512 3109 578 3119
rect 704 3109 770 3119
rect 896 3109 962 3119
rect 1088 3109 1154 3119
rect 1280 3109 1346 3119
rect 1472 3109 1528 3119
rect 1956 3109 2022 3119
rect 2148 3109 2214 3119
rect 2340 3109 2406 3119
rect 2532 3109 2598 3119
rect 2724 3109 2790 3119
rect 2916 3109 2982 3119
rect 3108 3109 3174 3119
rect 3300 3109 3356 3119
rect 3784 3109 3850 3119
rect 3976 3109 4042 3119
rect 4168 3109 4234 3119
rect 4360 3109 4426 3119
rect 4552 3109 4618 3119
rect 4744 3109 4810 3119
rect 4936 3109 5002 3119
rect 5128 3109 5184 3119
rect 5612 3109 5678 3119
rect 5804 3109 5870 3119
rect 5996 3109 6062 3119
rect 6188 3109 6254 3119
rect 6380 3109 6446 3119
rect 6572 3109 6638 3119
rect 6764 3109 6830 3119
rect 6956 3109 7012 3119
rect 7440 3109 7506 3119
rect 7632 3109 7698 3119
rect 7824 3109 7890 3119
rect 8016 3109 8082 3119
rect 8208 3109 8274 3119
rect 8400 3109 8466 3119
rect 8592 3109 8658 3119
rect 8784 3109 8840 3119
rect 9268 3109 9334 3119
rect 9460 3109 9526 3119
rect 9652 3109 9718 3119
rect 9844 3109 9910 3119
rect 10036 3109 10102 3119
rect 10228 3109 10294 3119
rect 10420 3109 10486 3119
rect 10612 3109 10668 3119
rect 11096 3109 11162 3119
rect 11288 3109 11354 3119
rect 11480 3109 11546 3119
rect 11672 3109 11738 3119
rect 11864 3109 11930 3119
rect 12056 3109 12122 3119
rect 12248 3109 12314 3119
rect 12440 3109 12496 3119
rect 12924 3109 12990 3119
rect 13116 3109 13182 3119
rect 13308 3109 13374 3119
rect 13500 3109 13566 3119
rect 13692 3109 13758 3119
rect 13884 3109 13950 3119
rect 14076 3109 14142 3119
rect 14268 3109 14324 3119
rect 14752 3109 14818 3119
rect 14944 3109 15010 3119
rect 15136 3109 15202 3119
rect 15328 3109 15394 3119
rect 15520 3109 15586 3119
rect 15712 3109 15778 3119
rect 15904 3109 15970 3119
rect 16096 3109 16152 3119
rect 16580 3109 16646 3119
rect 16772 3109 16838 3119
rect 16964 3109 17030 3119
rect 17156 3109 17222 3119
rect 17348 3109 17414 3119
rect 17540 3109 17606 3119
rect 17732 3109 17798 3119
rect 17924 3109 17980 3119
rect 18408 3109 18474 3119
rect 18600 3109 18666 3119
rect 18792 3109 18858 3119
rect 18984 3109 19050 3119
rect 19176 3109 19242 3119
rect 19368 3109 19434 3119
rect 19560 3109 19626 3119
rect 19752 3109 19808 3119
rect 20236 3109 20302 3119
rect 20428 3109 20494 3119
rect 20620 3109 20686 3119
rect 20812 3109 20878 3119
rect 21004 3109 21070 3119
rect 21196 3109 21262 3119
rect 21388 3109 21454 3119
rect 21580 3109 21636 3119
rect 0 2956 128 3109
rect 194 2956 320 3109
rect 386 2956 512 3109
rect 578 2956 704 3109
rect 770 2956 896 3109
rect 962 2956 1088 3109
rect 1154 2956 1280 3109
rect 1346 2956 1472 3109
rect 1528 2956 1708 3109
rect 1828 2956 1956 3109
rect 2022 2956 2148 3109
rect 2214 2956 2340 3109
rect 2406 2956 2532 3109
rect 2598 2956 2724 3109
rect 2790 2956 2916 3109
rect 2982 2956 3108 3109
rect 3174 2956 3300 3109
rect 3356 2956 3536 3109
rect 3656 2956 3784 3109
rect 3850 2956 3976 3109
rect 4042 2956 4168 3109
rect 4234 2956 4360 3109
rect 4426 2956 4552 3109
rect 4618 2956 4744 3109
rect 4810 2956 4936 3109
rect 5002 2956 5128 3109
rect 5184 2956 5364 3109
rect 5484 2956 5612 3109
rect 5678 2956 5804 3109
rect 5870 2956 5996 3109
rect 6062 2956 6188 3109
rect 6254 2956 6380 3109
rect 6446 2956 6572 3109
rect 6638 2956 6764 3109
rect 6830 2956 6956 3109
rect 7012 2956 7192 3109
rect 7312 2956 7440 3109
rect 7506 2956 7632 3109
rect 7698 2956 7824 3109
rect 7890 2956 8016 3109
rect 8082 2956 8208 3109
rect 8274 2956 8400 3109
rect 8466 2956 8592 3109
rect 8658 2956 8784 3109
rect 8840 2956 9020 3109
rect 9140 2956 9268 3109
rect 9334 2956 9460 3109
rect 9526 2956 9652 3109
rect 9718 2956 9844 3109
rect 9910 2956 10036 3109
rect 10102 2956 10228 3109
rect 10294 2956 10420 3109
rect 10486 2956 10612 3109
rect 10668 2956 10848 3109
rect 10968 2956 11096 3109
rect 11162 2956 11288 3109
rect 11354 2956 11480 3109
rect 11546 2956 11672 3109
rect 11738 2956 11864 3109
rect 11930 2956 12056 3109
rect 12122 2956 12248 3109
rect 12314 2956 12440 3109
rect 12496 2956 12676 3109
rect 12796 2956 12924 3109
rect 12990 2956 13116 3109
rect 13182 2956 13308 3109
rect 13374 2956 13500 3109
rect 13566 2956 13692 3109
rect 13758 2956 13884 3109
rect 13950 2956 14076 3109
rect 14142 2956 14268 3109
rect 14324 2956 14504 3109
rect 14624 2956 14752 3109
rect 14818 2956 14944 3109
rect 15010 2956 15136 3109
rect 15202 2956 15328 3109
rect 15394 2956 15520 3109
rect 15586 2956 15712 3109
rect 15778 2956 15904 3109
rect 15970 2956 16096 3109
rect 16152 2956 16332 3109
rect 16452 2956 16580 3109
rect 16646 2956 16772 3109
rect 16838 2956 16964 3109
rect 17030 2956 17156 3109
rect 17222 2956 17348 3109
rect 17414 2956 17540 3109
rect 17606 2956 17732 3109
rect 17798 2956 17924 3109
rect 17980 2956 18160 3109
rect 18280 2956 18408 3109
rect 18474 2956 18600 3109
rect 18666 2956 18792 3109
rect 18858 2956 18984 3109
rect 19050 2956 19176 3109
rect 19242 2956 19368 3109
rect 19434 2956 19560 3109
rect 19626 2956 19752 3109
rect 19808 2956 19988 3109
rect 20108 2956 20236 3109
rect 20302 2956 20428 3109
rect 20494 2956 20620 3109
rect 20686 2956 20812 3109
rect 20878 2956 21004 3109
rect 21070 2956 21196 3109
rect 21262 2956 21388 3109
rect 21454 2956 21580 3109
rect 21636 2956 21816 3109
rect 128 2946 194 2956
rect 320 2946 386 2956
rect 512 2946 578 2956
rect 704 2946 770 2956
rect 896 2946 962 2956
rect 1088 2946 1154 2956
rect 1280 2946 1346 2956
rect 1472 2946 1528 2956
rect 1956 2946 2022 2956
rect 2148 2946 2214 2956
rect 2340 2946 2406 2956
rect 2532 2946 2598 2956
rect 2724 2946 2790 2956
rect 2916 2946 2982 2956
rect 3108 2946 3174 2956
rect 3300 2946 3356 2956
rect 3784 2946 3850 2956
rect 3976 2946 4042 2956
rect 4168 2946 4234 2956
rect 4360 2946 4426 2956
rect 4552 2946 4618 2956
rect 4744 2946 4810 2956
rect 4936 2946 5002 2956
rect 5128 2946 5184 2956
rect 5612 2946 5678 2956
rect 5804 2946 5870 2956
rect 5996 2946 6062 2956
rect 6188 2946 6254 2956
rect 6380 2946 6446 2956
rect 6572 2946 6638 2956
rect 6764 2946 6830 2956
rect 6956 2946 7012 2956
rect 7440 2946 7506 2956
rect 7632 2946 7698 2956
rect 7824 2946 7890 2956
rect 8016 2946 8082 2956
rect 8208 2946 8274 2956
rect 8400 2946 8466 2956
rect 8592 2946 8658 2956
rect 8784 2946 8840 2956
rect 9268 2946 9334 2956
rect 9460 2946 9526 2956
rect 9652 2946 9718 2956
rect 9844 2946 9910 2956
rect 10036 2946 10102 2956
rect 10228 2946 10294 2956
rect 10420 2946 10486 2956
rect 10612 2946 10668 2956
rect 11096 2946 11162 2956
rect 11288 2946 11354 2956
rect 11480 2946 11546 2956
rect 11672 2946 11738 2956
rect 11864 2946 11930 2956
rect 12056 2946 12122 2956
rect 12248 2946 12314 2956
rect 12440 2946 12496 2956
rect 12924 2946 12990 2956
rect 13116 2946 13182 2956
rect 13308 2946 13374 2956
rect 13500 2946 13566 2956
rect 13692 2946 13758 2956
rect 13884 2946 13950 2956
rect 14076 2946 14142 2956
rect 14268 2946 14324 2956
rect 14752 2946 14818 2956
rect 14944 2946 15010 2956
rect 15136 2946 15202 2956
rect 15328 2946 15394 2956
rect 15520 2946 15586 2956
rect 15712 2946 15778 2956
rect 15904 2946 15970 2956
rect 16096 2946 16152 2956
rect 16580 2946 16646 2956
rect 16772 2946 16838 2956
rect 16964 2946 17030 2956
rect 17156 2946 17222 2956
rect 17348 2946 17414 2956
rect 17540 2946 17606 2956
rect 17732 2946 17798 2956
rect 17924 2946 17980 2956
rect 18408 2946 18474 2956
rect 18600 2946 18666 2956
rect 18792 2946 18858 2956
rect 18984 2946 19050 2956
rect 19176 2946 19242 2956
rect 19368 2946 19434 2956
rect 19560 2946 19626 2956
rect 19752 2946 19808 2956
rect 20236 2946 20302 2956
rect 20428 2946 20494 2956
rect 20620 2946 20686 2956
rect 20812 2946 20878 2956
rect 21004 2946 21070 2956
rect 21196 2946 21262 2956
rect 21388 2946 21454 2956
rect 21580 2946 21636 2956
rect 32 2608 98 2618
rect 224 2608 290 2618
rect 416 2608 482 2618
rect 608 2608 674 2618
rect 800 2608 866 2618
rect 992 2608 1058 2618
rect 1184 2608 1250 2618
rect 1376 2608 1442 2618
rect 1860 2608 1926 2618
rect 2052 2608 2118 2618
rect 2244 2608 2310 2618
rect 2436 2608 2502 2618
rect 2628 2608 2694 2618
rect 2820 2608 2886 2618
rect 3012 2608 3078 2618
rect 3204 2608 3270 2618
rect 3688 2608 3754 2618
rect 3880 2608 3946 2618
rect 4072 2608 4138 2618
rect 4264 2608 4330 2618
rect 4456 2608 4522 2618
rect 4648 2608 4714 2618
rect 4840 2608 4906 2618
rect 5032 2608 5098 2618
rect 5516 2608 5582 2618
rect 5708 2608 5774 2618
rect 5900 2608 5966 2618
rect 6092 2608 6158 2618
rect 6284 2608 6350 2618
rect 6476 2608 6542 2618
rect 6668 2608 6734 2618
rect 6860 2608 6926 2618
rect 7344 2608 7410 2618
rect 7536 2608 7602 2618
rect 7728 2608 7794 2618
rect 7920 2608 7986 2618
rect 8112 2608 8178 2618
rect 8304 2608 8370 2618
rect 8496 2608 8562 2618
rect 8688 2608 8754 2618
rect 9172 2608 9238 2618
rect 9364 2608 9430 2618
rect 9556 2608 9622 2618
rect 9748 2608 9814 2618
rect 9940 2608 10006 2618
rect 10132 2608 10198 2618
rect 10324 2608 10390 2618
rect 10516 2608 10582 2618
rect 11000 2608 11066 2618
rect 11192 2608 11258 2618
rect 11384 2608 11450 2618
rect 11576 2608 11642 2618
rect 11768 2608 11834 2618
rect 11960 2608 12026 2618
rect 12152 2608 12218 2618
rect 12344 2608 12410 2618
rect 12828 2608 12894 2618
rect 13020 2608 13086 2618
rect 13212 2608 13278 2618
rect 13404 2608 13470 2618
rect 13596 2608 13662 2618
rect 13788 2608 13854 2618
rect 13980 2608 14046 2618
rect 14172 2608 14238 2618
rect 14656 2608 14722 2618
rect 14848 2608 14914 2618
rect 15040 2608 15106 2618
rect 15232 2608 15298 2618
rect 15424 2608 15490 2618
rect 15616 2608 15682 2618
rect 15808 2608 15874 2618
rect 16000 2608 16066 2618
rect 16484 2608 16550 2618
rect 16676 2608 16742 2618
rect 16868 2608 16934 2618
rect 17060 2608 17126 2618
rect 17252 2608 17318 2618
rect 17444 2608 17510 2618
rect 17636 2608 17702 2618
rect 17828 2608 17894 2618
rect 18312 2608 18378 2618
rect 18504 2608 18570 2618
rect 18696 2608 18762 2618
rect 18888 2608 18954 2618
rect 19080 2608 19146 2618
rect 19272 2608 19338 2618
rect 19464 2608 19530 2618
rect 19656 2608 19722 2618
rect 20140 2608 20206 2618
rect 20332 2608 20398 2618
rect 20524 2608 20590 2618
rect 20716 2608 20782 2618
rect 20908 2608 20974 2618
rect 21100 2608 21166 2618
rect 21292 2608 21358 2618
rect 21484 2608 21550 2618
rect 0 2455 32 2608
rect 98 2455 224 2608
rect 290 2455 416 2608
rect 482 2455 608 2608
rect 674 2455 800 2608
rect 866 2455 992 2608
rect 1058 2455 1184 2608
rect 1250 2455 1376 2608
rect 1828 2455 1860 2608
rect 1926 2455 2052 2608
rect 2118 2455 2244 2608
rect 2310 2455 2436 2608
rect 2502 2455 2628 2608
rect 2694 2455 2820 2608
rect 2886 2455 3012 2608
rect 3078 2455 3204 2608
rect 3656 2455 3688 2608
rect 3754 2455 3880 2608
rect 3946 2455 4072 2608
rect 4138 2455 4264 2608
rect 4330 2455 4456 2608
rect 4522 2455 4648 2608
rect 4714 2455 4840 2608
rect 4906 2455 5032 2608
rect 5484 2455 5516 2608
rect 5582 2455 5708 2608
rect 5774 2455 5900 2608
rect 5966 2455 6092 2608
rect 6158 2455 6284 2608
rect 6350 2455 6476 2608
rect 6542 2455 6668 2608
rect 6734 2455 6860 2608
rect 7312 2455 7344 2608
rect 7410 2455 7536 2608
rect 7602 2455 7728 2608
rect 7794 2455 7920 2608
rect 7986 2455 8112 2608
rect 8178 2455 8304 2608
rect 8370 2455 8496 2608
rect 8562 2455 8688 2608
rect 9140 2455 9172 2608
rect 9238 2455 9364 2608
rect 9430 2455 9556 2608
rect 9622 2455 9748 2608
rect 9814 2455 9940 2608
rect 10006 2455 10132 2608
rect 10198 2455 10324 2608
rect 10390 2455 10516 2608
rect 10968 2455 11000 2608
rect 11066 2455 11192 2608
rect 11258 2455 11384 2608
rect 11450 2455 11576 2608
rect 11642 2455 11768 2608
rect 11834 2455 11960 2608
rect 12026 2455 12152 2608
rect 12218 2455 12344 2608
rect 12796 2455 12828 2608
rect 12894 2455 13020 2608
rect 13086 2455 13212 2608
rect 13278 2455 13404 2608
rect 13470 2455 13596 2608
rect 13662 2455 13788 2608
rect 13854 2455 13980 2608
rect 14046 2455 14172 2608
rect 14624 2455 14656 2608
rect 14722 2455 14848 2608
rect 14914 2455 15040 2608
rect 15106 2455 15232 2608
rect 15298 2455 15424 2608
rect 15490 2455 15616 2608
rect 15682 2455 15808 2608
rect 15874 2455 16000 2608
rect 16452 2455 16484 2608
rect 16550 2455 16676 2608
rect 16742 2455 16868 2608
rect 16934 2455 17060 2608
rect 17126 2455 17252 2608
rect 17318 2455 17444 2608
rect 17510 2455 17636 2608
rect 17702 2455 17828 2608
rect 18280 2455 18312 2608
rect 18378 2455 18504 2608
rect 18570 2455 18696 2608
rect 18762 2455 18888 2608
rect 18954 2455 19080 2608
rect 19146 2455 19272 2608
rect 19338 2455 19464 2608
rect 19530 2455 19656 2608
rect 20108 2455 20140 2608
rect 20206 2455 20332 2608
rect 20398 2455 20524 2608
rect 20590 2455 20716 2608
rect 20782 2455 20908 2608
rect 20974 2455 21100 2608
rect 21166 2455 21292 2608
rect 21358 2455 21484 2608
rect 32 2445 98 2455
rect 224 2445 290 2455
rect 416 2445 482 2455
rect 608 2445 674 2455
rect 800 2445 866 2455
rect 992 2445 1058 2455
rect 1184 2445 1250 2455
rect 1376 2445 1442 2455
rect 1860 2445 1926 2455
rect 2052 2445 2118 2455
rect 2244 2445 2310 2455
rect 2436 2445 2502 2455
rect 2628 2445 2694 2455
rect 2820 2445 2886 2455
rect 3012 2445 3078 2455
rect 3204 2445 3270 2455
rect 3688 2445 3754 2455
rect 3880 2445 3946 2455
rect 4072 2445 4138 2455
rect 4264 2445 4330 2455
rect 4456 2445 4522 2455
rect 4648 2445 4714 2455
rect 4840 2445 4906 2455
rect 5032 2445 5098 2455
rect 5516 2445 5582 2455
rect 5708 2445 5774 2455
rect 5900 2445 5966 2455
rect 6092 2445 6158 2455
rect 6284 2445 6350 2455
rect 6476 2445 6542 2455
rect 6668 2445 6734 2455
rect 6860 2445 6926 2455
rect 7344 2445 7410 2455
rect 7536 2445 7602 2455
rect 7728 2445 7794 2455
rect 7920 2445 7986 2455
rect 8112 2445 8178 2455
rect 8304 2445 8370 2455
rect 8496 2445 8562 2455
rect 8688 2445 8754 2455
rect 9172 2445 9238 2455
rect 9364 2445 9430 2455
rect 9556 2445 9622 2455
rect 9748 2445 9814 2455
rect 9940 2445 10006 2455
rect 10132 2445 10198 2455
rect 10324 2445 10390 2455
rect 10516 2445 10582 2455
rect 11000 2445 11066 2455
rect 11192 2445 11258 2455
rect 11384 2445 11450 2455
rect 11576 2445 11642 2455
rect 11768 2445 11834 2455
rect 11960 2445 12026 2455
rect 12152 2445 12218 2455
rect 12344 2445 12410 2455
rect 12828 2445 12894 2455
rect 13020 2445 13086 2455
rect 13212 2445 13278 2455
rect 13404 2445 13470 2455
rect 13596 2445 13662 2455
rect 13788 2445 13854 2455
rect 13980 2445 14046 2455
rect 14172 2445 14238 2455
rect 14656 2445 14722 2455
rect 14848 2445 14914 2455
rect 15040 2445 15106 2455
rect 15232 2445 15298 2455
rect 15424 2445 15490 2455
rect 15616 2445 15682 2455
rect 15808 2445 15874 2455
rect 16000 2445 16066 2455
rect 16484 2445 16550 2455
rect 16676 2445 16742 2455
rect 16868 2445 16934 2455
rect 17060 2445 17126 2455
rect 17252 2445 17318 2455
rect 17444 2445 17510 2455
rect 17636 2445 17702 2455
rect 17828 2445 17894 2455
rect 18312 2445 18378 2455
rect 18504 2445 18570 2455
rect 18696 2445 18762 2455
rect 18888 2445 18954 2455
rect 19080 2445 19146 2455
rect 19272 2445 19338 2455
rect 19464 2445 19530 2455
rect 19656 2445 19722 2455
rect 20140 2445 20206 2455
rect 20332 2445 20398 2455
rect 20524 2445 20590 2455
rect 20716 2445 20782 2455
rect 20908 2445 20974 2455
rect 21100 2445 21166 2455
rect 21292 2445 21358 2455
rect 21484 2445 21550 2455
rect 128 2395 194 2405
rect 320 2395 386 2405
rect 512 2395 578 2405
rect 704 2395 770 2405
rect 896 2395 962 2405
rect 1088 2395 1154 2405
rect 1280 2395 1346 2405
rect 1472 2395 1528 2405
rect 1956 2395 2022 2405
rect 2148 2395 2214 2405
rect 2340 2395 2406 2405
rect 2532 2395 2598 2405
rect 2724 2395 2790 2405
rect 2916 2395 2982 2405
rect 3108 2395 3174 2405
rect 3300 2395 3356 2405
rect 3784 2395 3850 2405
rect 3976 2395 4042 2405
rect 4168 2395 4234 2405
rect 4360 2395 4426 2405
rect 4552 2395 4618 2405
rect 4744 2395 4810 2405
rect 4936 2395 5002 2405
rect 5128 2395 5184 2405
rect 5612 2395 5678 2405
rect 5804 2395 5870 2405
rect 5996 2395 6062 2405
rect 6188 2395 6254 2405
rect 6380 2395 6446 2405
rect 6572 2395 6638 2405
rect 6764 2395 6830 2405
rect 6956 2395 7012 2405
rect 7440 2395 7506 2405
rect 7632 2395 7698 2405
rect 7824 2395 7890 2405
rect 8016 2395 8082 2405
rect 8208 2395 8274 2405
rect 8400 2395 8466 2405
rect 8592 2395 8658 2405
rect 8784 2395 8840 2405
rect 9268 2395 9334 2405
rect 9460 2395 9526 2405
rect 9652 2395 9718 2405
rect 9844 2395 9910 2405
rect 10036 2395 10102 2405
rect 10228 2395 10294 2405
rect 10420 2395 10486 2405
rect 10612 2395 10668 2405
rect 11096 2395 11162 2405
rect 11288 2395 11354 2405
rect 11480 2395 11546 2405
rect 11672 2395 11738 2405
rect 11864 2395 11930 2405
rect 12056 2395 12122 2405
rect 12248 2395 12314 2405
rect 12440 2395 12496 2405
rect 12924 2395 12990 2405
rect 13116 2395 13182 2405
rect 13308 2395 13374 2405
rect 13500 2395 13566 2405
rect 13692 2395 13758 2405
rect 13884 2395 13950 2405
rect 14076 2395 14142 2405
rect 14268 2395 14324 2405
rect 14752 2395 14818 2405
rect 14944 2395 15010 2405
rect 15136 2395 15202 2405
rect 15328 2395 15394 2405
rect 15520 2395 15586 2405
rect 15712 2395 15778 2405
rect 15904 2395 15970 2405
rect 16096 2395 16152 2405
rect 16580 2395 16646 2405
rect 16772 2395 16838 2405
rect 16964 2395 17030 2405
rect 17156 2395 17222 2405
rect 17348 2395 17414 2405
rect 17540 2395 17606 2405
rect 17732 2395 17798 2405
rect 17924 2395 17980 2405
rect 18408 2395 18474 2405
rect 18600 2395 18666 2405
rect 18792 2395 18858 2405
rect 18984 2395 19050 2405
rect 19176 2395 19242 2405
rect 19368 2395 19434 2405
rect 19560 2395 19626 2405
rect 19752 2395 19808 2405
rect 20236 2395 20302 2405
rect 20428 2395 20494 2405
rect 20620 2395 20686 2405
rect 20812 2395 20878 2405
rect 21004 2395 21070 2405
rect 21196 2395 21262 2405
rect 21388 2395 21454 2405
rect 21580 2395 21636 2405
rect 0 2242 128 2395
rect 194 2242 320 2395
rect 386 2242 512 2395
rect 578 2242 704 2395
rect 770 2242 896 2395
rect 962 2242 1088 2395
rect 1154 2242 1280 2395
rect 1346 2242 1472 2395
rect 1528 2242 1708 2395
rect 1828 2242 1956 2395
rect 2022 2242 2148 2395
rect 2214 2242 2340 2395
rect 2406 2242 2532 2395
rect 2598 2242 2724 2395
rect 2790 2242 2916 2395
rect 2982 2242 3108 2395
rect 3174 2242 3300 2395
rect 3356 2242 3536 2395
rect 3656 2242 3784 2395
rect 3850 2242 3976 2395
rect 4042 2242 4168 2395
rect 4234 2242 4360 2395
rect 4426 2242 4552 2395
rect 4618 2242 4744 2395
rect 4810 2242 4936 2395
rect 5002 2242 5128 2395
rect 5184 2242 5364 2395
rect 5484 2242 5612 2395
rect 5678 2242 5804 2395
rect 5870 2242 5996 2395
rect 6062 2242 6188 2395
rect 6254 2242 6380 2395
rect 6446 2242 6572 2395
rect 6638 2242 6764 2395
rect 6830 2242 6956 2395
rect 7012 2242 7192 2395
rect 7312 2242 7440 2395
rect 7506 2242 7632 2395
rect 7698 2242 7824 2395
rect 7890 2242 8016 2395
rect 8082 2242 8208 2395
rect 8274 2242 8400 2395
rect 8466 2242 8592 2395
rect 8658 2242 8784 2395
rect 8840 2242 9020 2395
rect 9140 2242 9268 2395
rect 9334 2242 9460 2395
rect 9526 2242 9652 2395
rect 9718 2242 9844 2395
rect 9910 2242 10036 2395
rect 10102 2242 10228 2395
rect 10294 2242 10420 2395
rect 10486 2242 10612 2395
rect 10668 2242 10848 2395
rect 10968 2242 11096 2395
rect 11162 2242 11288 2395
rect 11354 2242 11480 2395
rect 11546 2242 11672 2395
rect 11738 2242 11864 2395
rect 11930 2242 12056 2395
rect 12122 2242 12248 2395
rect 12314 2242 12440 2395
rect 12496 2242 12676 2395
rect 12796 2242 12924 2395
rect 12990 2242 13116 2395
rect 13182 2242 13308 2395
rect 13374 2242 13500 2395
rect 13566 2242 13692 2395
rect 13758 2242 13884 2395
rect 13950 2242 14076 2395
rect 14142 2242 14268 2395
rect 14324 2242 14504 2395
rect 14624 2242 14752 2395
rect 14818 2242 14944 2395
rect 15010 2242 15136 2395
rect 15202 2242 15328 2395
rect 15394 2242 15520 2395
rect 15586 2242 15712 2395
rect 15778 2242 15904 2395
rect 15970 2242 16096 2395
rect 16152 2242 16332 2395
rect 16452 2242 16580 2395
rect 16646 2242 16772 2395
rect 16838 2242 16964 2395
rect 17030 2242 17156 2395
rect 17222 2242 17348 2395
rect 17414 2242 17540 2395
rect 17606 2242 17732 2395
rect 17798 2242 17924 2395
rect 17980 2242 18160 2395
rect 18280 2242 18408 2395
rect 18474 2242 18600 2395
rect 18666 2242 18792 2395
rect 18858 2242 18984 2395
rect 19050 2242 19176 2395
rect 19242 2242 19368 2395
rect 19434 2242 19560 2395
rect 19626 2242 19752 2395
rect 19808 2242 19988 2395
rect 20108 2242 20236 2395
rect 20302 2242 20428 2395
rect 20494 2242 20620 2395
rect 20686 2242 20812 2395
rect 20878 2242 21004 2395
rect 21070 2242 21196 2395
rect 21262 2242 21388 2395
rect 21454 2242 21580 2395
rect 21636 2242 21816 2395
rect 128 2232 194 2242
rect 320 2232 386 2242
rect 512 2232 578 2242
rect 704 2232 770 2242
rect 896 2232 962 2242
rect 1088 2232 1154 2242
rect 1280 2232 1346 2242
rect 1472 2232 1528 2242
rect 1956 2232 2022 2242
rect 2148 2232 2214 2242
rect 2340 2232 2406 2242
rect 2532 2232 2598 2242
rect 2724 2232 2790 2242
rect 2916 2232 2982 2242
rect 3108 2232 3174 2242
rect 3300 2232 3356 2242
rect 3784 2232 3850 2242
rect 3976 2232 4042 2242
rect 4168 2232 4234 2242
rect 4360 2232 4426 2242
rect 4552 2232 4618 2242
rect 4744 2232 4810 2242
rect 4936 2232 5002 2242
rect 5128 2232 5184 2242
rect 5612 2232 5678 2242
rect 5804 2232 5870 2242
rect 5996 2232 6062 2242
rect 6188 2232 6254 2242
rect 6380 2232 6446 2242
rect 6572 2232 6638 2242
rect 6764 2232 6830 2242
rect 6956 2232 7012 2242
rect 7440 2232 7506 2242
rect 7632 2232 7698 2242
rect 7824 2232 7890 2242
rect 8016 2232 8082 2242
rect 8208 2232 8274 2242
rect 8400 2232 8466 2242
rect 8592 2232 8658 2242
rect 8784 2232 8840 2242
rect 9268 2232 9334 2242
rect 9460 2232 9526 2242
rect 9652 2232 9718 2242
rect 9844 2232 9910 2242
rect 10036 2232 10102 2242
rect 10228 2232 10294 2242
rect 10420 2232 10486 2242
rect 10612 2232 10668 2242
rect 11096 2232 11162 2242
rect 11288 2232 11354 2242
rect 11480 2232 11546 2242
rect 11672 2232 11738 2242
rect 11864 2232 11930 2242
rect 12056 2232 12122 2242
rect 12248 2232 12314 2242
rect 12440 2232 12496 2242
rect 12924 2232 12990 2242
rect 13116 2232 13182 2242
rect 13308 2232 13374 2242
rect 13500 2232 13566 2242
rect 13692 2232 13758 2242
rect 13884 2232 13950 2242
rect 14076 2232 14142 2242
rect 14268 2232 14324 2242
rect 14752 2232 14818 2242
rect 14944 2232 15010 2242
rect 15136 2232 15202 2242
rect 15328 2232 15394 2242
rect 15520 2232 15586 2242
rect 15712 2232 15778 2242
rect 15904 2232 15970 2242
rect 16096 2232 16152 2242
rect 16580 2232 16646 2242
rect 16772 2232 16838 2242
rect 16964 2232 17030 2242
rect 17156 2232 17222 2242
rect 17348 2232 17414 2242
rect 17540 2232 17606 2242
rect 17732 2232 17798 2242
rect 17924 2232 17980 2242
rect 18408 2232 18474 2242
rect 18600 2232 18666 2242
rect 18792 2232 18858 2242
rect 18984 2232 19050 2242
rect 19176 2232 19242 2242
rect 19368 2232 19434 2242
rect 19560 2232 19626 2242
rect 19752 2232 19808 2242
rect 20236 2232 20302 2242
rect 20428 2232 20494 2242
rect 20620 2232 20686 2242
rect 20812 2232 20878 2242
rect 21004 2232 21070 2242
rect 21196 2232 21262 2242
rect 21388 2232 21454 2242
rect 21580 2232 21636 2242
rect 32 1894 98 1904
rect 224 1894 290 1904
rect 416 1894 482 1904
rect 608 1894 674 1904
rect 800 1894 866 1904
rect 992 1894 1058 1904
rect 1184 1894 1250 1904
rect 1376 1894 1442 1904
rect 1860 1894 1926 1904
rect 2052 1894 2118 1904
rect 2244 1894 2310 1904
rect 2436 1894 2502 1904
rect 2628 1894 2694 1904
rect 2820 1894 2886 1904
rect 3012 1894 3078 1904
rect 3204 1894 3270 1904
rect 3688 1894 3754 1904
rect 3880 1894 3946 1904
rect 4072 1894 4138 1904
rect 4264 1894 4330 1904
rect 4456 1894 4522 1904
rect 4648 1894 4714 1904
rect 4840 1894 4906 1904
rect 5032 1894 5098 1904
rect 5516 1894 5582 1904
rect 5708 1894 5774 1904
rect 5900 1894 5966 1904
rect 6092 1894 6158 1904
rect 6284 1894 6350 1904
rect 6476 1894 6542 1904
rect 6668 1894 6734 1904
rect 6860 1894 6926 1904
rect 7344 1894 7410 1904
rect 7536 1894 7602 1904
rect 7728 1894 7794 1904
rect 7920 1894 7986 1904
rect 8112 1894 8178 1904
rect 8304 1894 8370 1904
rect 8496 1894 8562 1904
rect 8688 1894 8754 1904
rect 9172 1894 9238 1904
rect 9364 1894 9430 1904
rect 9556 1894 9622 1904
rect 9748 1894 9814 1904
rect 9940 1894 10006 1904
rect 10132 1894 10198 1904
rect 10324 1894 10390 1904
rect 10516 1894 10582 1904
rect 11000 1894 11066 1904
rect 11192 1894 11258 1904
rect 11384 1894 11450 1904
rect 11576 1894 11642 1904
rect 11768 1894 11834 1904
rect 11960 1894 12026 1904
rect 12152 1894 12218 1904
rect 12344 1894 12410 1904
rect 12828 1894 12894 1904
rect 13020 1894 13086 1904
rect 13212 1894 13278 1904
rect 13404 1894 13470 1904
rect 13596 1894 13662 1904
rect 13788 1894 13854 1904
rect 13980 1894 14046 1904
rect 14172 1894 14238 1904
rect 14656 1894 14722 1904
rect 14848 1894 14914 1904
rect 15040 1894 15106 1904
rect 15232 1894 15298 1904
rect 15424 1894 15490 1904
rect 15616 1894 15682 1904
rect 15808 1894 15874 1904
rect 16000 1894 16066 1904
rect 16484 1894 16550 1904
rect 16676 1894 16742 1904
rect 16868 1894 16934 1904
rect 17060 1894 17126 1904
rect 17252 1894 17318 1904
rect 17444 1894 17510 1904
rect 17636 1894 17702 1904
rect 17828 1894 17894 1904
rect 18312 1894 18378 1904
rect 18504 1894 18570 1904
rect 18696 1894 18762 1904
rect 18888 1894 18954 1904
rect 19080 1894 19146 1904
rect 19272 1894 19338 1904
rect 19464 1894 19530 1904
rect 19656 1894 19722 1904
rect 20140 1894 20206 1904
rect 20332 1894 20398 1904
rect 20524 1894 20590 1904
rect 20716 1894 20782 1904
rect 20908 1894 20974 1904
rect 21100 1894 21166 1904
rect 21292 1894 21358 1904
rect 21484 1894 21550 1904
rect 0 1741 32 1894
rect 98 1741 224 1894
rect 290 1741 416 1894
rect 482 1741 608 1894
rect 674 1741 800 1894
rect 866 1741 992 1894
rect 1058 1741 1184 1894
rect 1250 1741 1376 1894
rect 1828 1741 1860 1894
rect 1926 1741 2052 1894
rect 2118 1741 2244 1894
rect 2310 1741 2436 1894
rect 2502 1741 2628 1894
rect 2694 1741 2820 1894
rect 2886 1741 3012 1894
rect 3078 1741 3204 1894
rect 3656 1741 3688 1894
rect 3754 1741 3880 1894
rect 3946 1741 4072 1894
rect 4138 1741 4264 1894
rect 4330 1741 4456 1894
rect 4522 1741 4648 1894
rect 4714 1741 4840 1894
rect 4906 1741 5032 1894
rect 5484 1741 5516 1894
rect 5582 1741 5708 1894
rect 5774 1741 5900 1894
rect 5966 1741 6092 1894
rect 6158 1741 6284 1894
rect 6350 1741 6476 1894
rect 6542 1741 6668 1894
rect 6734 1741 6860 1894
rect 7312 1741 7344 1894
rect 7410 1741 7536 1894
rect 7602 1741 7728 1894
rect 7794 1741 7920 1894
rect 7986 1741 8112 1894
rect 8178 1741 8304 1894
rect 8370 1741 8496 1894
rect 8562 1741 8688 1894
rect 9140 1741 9172 1894
rect 9238 1741 9364 1894
rect 9430 1741 9556 1894
rect 9622 1741 9748 1894
rect 9814 1741 9940 1894
rect 10006 1741 10132 1894
rect 10198 1741 10324 1894
rect 10390 1741 10516 1894
rect 10968 1741 11000 1894
rect 11066 1741 11192 1894
rect 11258 1741 11384 1894
rect 11450 1741 11576 1894
rect 11642 1741 11768 1894
rect 11834 1741 11960 1894
rect 12026 1741 12152 1894
rect 12218 1741 12344 1894
rect 12796 1741 12828 1894
rect 12894 1741 13020 1894
rect 13086 1741 13212 1894
rect 13278 1741 13404 1894
rect 13470 1741 13596 1894
rect 13662 1741 13788 1894
rect 13854 1741 13980 1894
rect 14046 1741 14172 1894
rect 14624 1741 14656 1894
rect 14722 1741 14848 1894
rect 14914 1741 15040 1894
rect 15106 1741 15232 1894
rect 15298 1741 15424 1894
rect 15490 1741 15616 1894
rect 15682 1741 15808 1894
rect 15874 1741 16000 1894
rect 16452 1741 16484 1894
rect 16550 1741 16676 1894
rect 16742 1741 16868 1894
rect 16934 1741 17060 1894
rect 17126 1741 17252 1894
rect 17318 1741 17444 1894
rect 17510 1741 17636 1894
rect 17702 1741 17828 1894
rect 18280 1741 18312 1894
rect 18378 1741 18504 1894
rect 18570 1741 18696 1894
rect 18762 1741 18888 1894
rect 18954 1741 19080 1894
rect 19146 1741 19272 1894
rect 19338 1741 19464 1894
rect 19530 1741 19656 1894
rect 20108 1741 20140 1894
rect 20206 1741 20332 1894
rect 20398 1741 20524 1894
rect 20590 1741 20716 1894
rect 20782 1741 20908 1894
rect 20974 1741 21100 1894
rect 21166 1741 21292 1894
rect 21358 1741 21484 1894
rect 32 1731 98 1741
rect 224 1731 290 1741
rect 416 1731 482 1741
rect 608 1731 674 1741
rect 800 1731 866 1741
rect 992 1731 1058 1741
rect 1184 1731 1250 1741
rect 1376 1731 1442 1741
rect 1860 1731 1926 1741
rect 2052 1731 2118 1741
rect 2244 1731 2310 1741
rect 2436 1731 2502 1741
rect 2628 1731 2694 1741
rect 2820 1731 2886 1741
rect 3012 1731 3078 1741
rect 3204 1731 3270 1741
rect 3688 1731 3754 1741
rect 3880 1731 3946 1741
rect 4072 1731 4138 1741
rect 4264 1731 4330 1741
rect 4456 1731 4522 1741
rect 4648 1731 4714 1741
rect 4840 1731 4906 1741
rect 5032 1731 5098 1741
rect 5516 1731 5582 1741
rect 5708 1731 5774 1741
rect 5900 1731 5966 1741
rect 6092 1731 6158 1741
rect 6284 1731 6350 1741
rect 6476 1731 6542 1741
rect 6668 1731 6734 1741
rect 6860 1731 6926 1741
rect 7344 1731 7410 1741
rect 7536 1731 7602 1741
rect 7728 1731 7794 1741
rect 7920 1731 7986 1741
rect 8112 1731 8178 1741
rect 8304 1731 8370 1741
rect 8496 1731 8562 1741
rect 8688 1731 8754 1741
rect 9172 1731 9238 1741
rect 9364 1731 9430 1741
rect 9556 1731 9622 1741
rect 9748 1731 9814 1741
rect 9940 1731 10006 1741
rect 10132 1731 10198 1741
rect 10324 1731 10390 1741
rect 10516 1731 10582 1741
rect 11000 1731 11066 1741
rect 11192 1731 11258 1741
rect 11384 1731 11450 1741
rect 11576 1731 11642 1741
rect 11768 1731 11834 1741
rect 11960 1731 12026 1741
rect 12152 1731 12218 1741
rect 12344 1731 12410 1741
rect 12828 1731 12894 1741
rect 13020 1731 13086 1741
rect 13212 1731 13278 1741
rect 13404 1731 13470 1741
rect 13596 1731 13662 1741
rect 13788 1731 13854 1741
rect 13980 1731 14046 1741
rect 14172 1731 14238 1741
rect 14656 1731 14722 1741
rect 14848 1731 14914 1741
rect 15040 1731 15106 1741
rect 15232 1731 15298 1741
rect 15424 1731 15490 1741
rect 15616 1731 15682 1741
rect 15808 1731 15874 1741
rect 16000 1731 16066 1741
rect 16484 1731 16550 1741
rect 16676 1731 16742 1741
rect 16868 1731 16934 1741
rect 17060 1731 17126 1741
rect 17252 1731 17318 1741
rect 17444 1731 17510 1741
rect 17636 1731 17702 1741
rect 17828 1731 17894 1741
rect 18312 1731 18378 1741
rect 18504 1731 18570 1741
rect 18696 1731 18762 1741
rect 18888 1731 18954 1741
rect 19080 1731 19146 1741
rect 19272 1731 19338 1741
rect 19464 1731 19530 1741
rect 19656 1731 19722 1741
rect 20140 1731 20206 1741
rect 20332 1731 20398 1741
rect 20524 1731 20590 1741
rect 20716 1731 20782 1741
rect 20908 1731 20974 1741
rect 21100 1731 21166 1741
rect 21292 1731 21358 1741
rect 21484 1731 21550 1741
rect 128 1681 194 1691
rect 320 1681 386 1691
rect 512 1681 578 1691
rect 704 1681 770 1691
rect 896 1681 962 1691
rect 1088 1681 1154 1691
rect 1280 1681 1346 1691
rect 1472 1681 1528 1691
rect 1956 1681 2022 1691
rect 2148 1681 2214 1691
rect 2340 1681 2406 1691
rect 2532 1681 2598 1691
rect 2724 1681 2790 1691
rect 2916 1681 2982 1691
rect 3108 1681 3174 1691
rect 3300 1681 3356 1691
rect 3784 1681 3850 1691
rect 3976 1681 4042 1691
rect 4168 1681 4234 1691
rect 4360 1681 4426 1691
rect 4552 1681 4618 1691
rect 4744 1681 4810 1691
rect 4936 1681 5002 1691
rect 5128 1681 5184 1691
rect 5612 1681 5678 1691
rect 5804 1681 5870 1691
rect 5996 1681 6062 1691
rect 6188 1681 6254 1691
rect 6380 1681 6446 1691
rect 6572 1681 6638 1691
rect 6764 1681 6830 1691
rect 6956 1681 7012 1691
rect 7440 1681 7506 1691
rect 7632 1681 7698 1691
rect 7824 1681 7890 1691
rect 8016 1681 8082 1691
rect 8208 1681 8274 1691
rect 8400 1681 8466 1691
rect 8592 1681 8658 1691
rect 8784 1681 8840 1691
rect 9268 1681 9334 1691
rect 9460 1681 9526 1691
rect 9652 1681 9718 1691
rect 9844 1681 9910 1691
rect 10036 1681 10102 1691
rect 10228 1681 10294 1691
rect 10420 1681 10486 1691
rect 10612 1681 10668 1691
rect 11096 1681 11162 1691
rect 11288 1681 11354 1691
rect 11480 1681 11546 1691
rect 11672 1681 11738 1691
rect 11864 1681 11930 1691
rect 12056 1681 12122 1691
rect 12248 1681 12314 1691
rect 12440 1681 12496 1691
rect 12924 1681 12990 1691
rect 13116 1681 13182 1691
rect 13308 1681 13374 1691
rect 13500 1681 13566 1691
rect 13692 1681 13758 1691
rect 13884 1681 13950 1691
rect 14076 1681 14142 1691
rect 14268 1681 14324 1691
rect 14752 1681 14818 1691
rect 14944 1681 15010 1691
rect 15136 1681 15202 1691
rect 15328 1681 15394 1691
rect 15520 1681 15586 1691
rect 15712 1681 15778 1691
rect 15904 1681 15970 1691
rect 16096 1681 16152 1691
rect 16580 1681 16646 1691
rect 16772 1681 16838 1691
rect 16964 1681 17030 1691
rect 17156 1681 17222 1691
rect 17348 1681 17414 1691
rect 17540 1681 17606 1691
rect 17732 1681 17798 1691
rect 17924 1681 17980 1691
rect 18408 1681 18474 1691
rect 18600 1681 18666 1691
rect 18792 1681 18858 1691
rect 18984 1681 19050 1691
rect 19176 1681 19242 1691
rect 19368 1681 19434 1691
rect 19560 1681 19626 1691
rect 19752 1681 19808 1691
rect 20236 1681 20302 1691
rect 20428 1681 20494 1691
rect 20620 1681 20686 1691
rect 20812 1681 20878 1691
rect 21004 1681 21070 1691
rect 21196 1681 21262 1691
rect 21388 1681 21454 1691
rect 21580 1681 21636 1691
rect 0 1528 128 1681
rect 194 1528 320 1681
rect 386 1528 512 1681
rect 578 1528 704 1681
rect 770 1528 896 1681
rect 962 1528 1088 1681
rect 1154 1528 1280 1681
rect 1346 1528 1472 1681
rect 1528 1528 1708 1681
rect 1828 1528 1956 1681
rect 2022 1528 2148 1681
rect 2214 1528 2340 1681
rect 2406 1528 2532 1681
rect 2598 1528 2724 1681
rect 2790 1528 2916 1681
rect 2982 1528 3108 1681
rect 3174 1528 3300 1681
rect 3356 1528 3536 1681
rect 3656 1528 3784 1681
rect 3850 1528 3976 1681
rect 4042 1528 4168 1681
rect 4234 1528 4360 1681
rect 4426 1528 4552 1681
rect 4618 1528 4744 1681
rect 4810 1528 4936 1681
rect 5002 1528 5128 1681
rect 5184 1528 5364 1681
rect 5484 1528 5612 1681
rect 5678 1528 5804 1681
rect 5870 1528 5996 1681
rect 6062 1528 6188 1681
rect 6254 1528 6380 1681
rect 6446 1528 6572 1681
rect 6638 1528 6764 1681
rect 6830 1528 6956 1681
rect 7012 1528 7192 1681
rect 7312 1528 7440 1681
rect 7506 1528 7632 1681
rect 7698 1528 7824 1681
rect 7890 1528 8016 1681
rect 8082 1528 8208 1681
rect 8274 1528 8400 1681
rect 8466 1528 8592 1681
rect 8658 1528 8784 1681
rect 8840 1528 9020 1681
rect 9140 1528 9268 1681
rect 9334 1528 9460 1681
rect 9526 1528 9652 1681
rect 9718 1528 9844 1681
rect 9910 1528 10036 1681
rect 10102 1528 10228 1681
rect 10294 1528 10420 1681
rect 10486 1528 10612 1681
rect 10668 1528 10848 1681
rect 10968 1528 11096 1681
rect 11162 1528 11288 1681
rect 11354 1528 11480 1681
rect 11546 1528 11672 1681
rect 11738 1528 11864 1681
rect 11930 1528 12056 1681
rect 12122 1528 12248 1681
rect 12314 1528 12440 1681
rect 12496 1528 12676 1681
rect 12796 1528 12924 1681
rect 12990 1528 13116 1681
rect 13182 1528 13308 1681
rect 13374 1528 13500 1681
rect 13566 1528 13692 1681
rect 13758 1528 13884 1681
rect 13950 1528 14076 1681
rect 14142 1528 14268 1681
rect 14324 1528 14504 1681
rect 14624 1528 14752 1681
rect 14818 1528 14944 1681
rect 15010 1528 15136 1681
rect 15202 1528 15328 1681
rect 15394 1528 15520 1681
rect 15586 1528 15712 1681
rect 15778 1528 15904 1681
rect 15970 1528 16096 1681
rect 16152 1528 16332 1681
rect 16452 1528 16580 1681
rect 16646 1528 16772 1681
rect 16838 1528 16964 1681
rect 17030 1528 17156 1681
rect 17222 1528 17348 1681
rect 17414 1528 17540 1681
rect 17606 1528 17732 1681
rect 17798 1528 17924 1681
rect 17980 1528 18160 1681
rect 18280 1528 18408 1681
rect 18474 1528 18600 1681
rect 18666 1528 18792 1681
rect 18858 1528 18984 1681
rect 19050 1528 19176 1681
rect 19242 1528 19368 1681
rect 19434 1528 19560 1681
rect 19626 1528 19752 1681
rect 19808 1528 19988 1681
rect 20108 1528 20236 1681
rect 20302 1528 20428 1681
rect 20494 1528 20620 1681
rect 20686 1528 20812 1681
rect 20878 1528 21004 1681
rect 21070 1528 21196 1681
rect 21262 1528 21388 1681
rect 21454 1528 21580 1681
rect 21636 1528 21816 1681
rect 128 1518 194 1528
rect 320 1518 386 1528
rect 512 1518 578 1528
rect 704 1518 770 1528
rect 896 1518 962 1528
rect 1088 1518 1154 1528
rect 1280 1518 1346 1528
rect 1472 1518 1528 1528
rect 1956 1518 2022 1528
rect 2148 1518 2214 1528
rect 2340 1518 2406 1528
rect 2532 1518 2598 1528
rect 2724 1518 2790 1528
rect 2916 1518 2982 1528
rect 3108 1518 3174 1528
rect 3300 1518 3356 1528
rect 3784 1518 3850 1528
rect 3976 1518 4042 1528
rect 4168 1518 4234 1528
rect 4360 1518 4426 1528
rect 4552 1518 4618 1528
rect 4744 1518 4810 1528
rect 4936 1518 5002 1528
rect 5128 1518 5184 1528
rect 5612 1518 5678 1528
rect 5804 1518 5870 1528
rect 5996 1518 6062 1528
rect 6188 1518 6254 1528
rect 6380 1518 6446 1528
rect 6572 1518 6638 1528
rect 6764 1518 6830 1528
rect 6956 1518 7012 1528
rect 7440 1518 7506 1528
rect 7632 1518 7698 1528
rect 7824 1518 7890 1528
rect 8016 1518 8082 1528
rect 8208 1518 8274 1528
rect 8400 1518 8466 1528
rect 8592 1518 8658 1528
rect 8784 1518 8840 1528
rect 9268 1518 9334 1528
rect 9460 1518 9526 1528
rect 9652 1518 9718 1528
rect 9844 1518 9910 1528
rect 10036 1518 10102 1528
rect 10228 1518 10294 1528
rect 10420 1518 10486 1528
rect 10612 1518 10668 1528
rect 11096 1518 11162 1528
rect 11288 1518 11354 1528
rect 11480 1518 11546 1528
rect 11672 1518 11738 1528
rect 11864 1518 11930 1528
rect 12056 1518 12122 1528
rect 12248 1518 12314 1528
rect 12440 1518 12496 1528
rect 12924 1518 12990 1528
rect 13116 1518 13182 1528
rect 13308 1518 13374 1528
rect 13500 1518 13566 1528
rect 13692 1518 13758 1528
rect 13884 1518 13950 1528
rect 14076 1518 14142 1528
rect 14268 1518 14324 1528
rect 14752 1518 14818 1528
rect 14944 1518 15010 1528
rect 15136 1518 15202 1528
rect 15328 1518 15394 1528
rect 15520 1518 15586 1528
rect 15712 1518 15778 1528
rect 15904 1518 15970 1528
rect 16096 1518 16152 1528
rect 16580 1518 16646 1528
rect 16772 1518 16838 1528
rect 16964 1518 17030 1528
rect 17156 1518 17222 1528
rect 17348 1518 17414 1528
rect 17540 1518 17606 1528
rect 17732 1518 17798 1528
rect 17924 1518 17980 1528
rect 18408 1518 18474 1528
rect 18600 1518 18666 1528
rect 18792 1518 18858 1528
rect 18984 1518 19050 1528
rect 19176 1518 19242 1528
rect 19368 1518 19434 1528
rect 19560 1518 19626 1528
rect 19752 1518 19808 1528
rect 20236 1518 20302 1528
rect 20428 1518 20494 1528
rect 20620 1518 20686 1528
rect 20812 1518 20878 1528
rect 21004 1518 21070 1528
rect 21196 1518 21262 1528
rect 21388 1518 21454 1528
rect 21580 1518 21636 1528
rect 32 1180 98 1190
rect 224 1180 290 1190
rect 416 1180 482 1190
rect 608 1180 674 1190
rect 800 1180 866 1190
rect 992 1180 1058 1190
rect 1184 1180 1250 1190
rect 1376 1180 1442 1190
rect 1860 1180 1926 1190
rect 2052 1180 2118 1190
rect 2244 1180 2310 1190
rect 2436 1180 2502 1190
rect 2628 1180 2694 1190
rect 2820 1180 2886 1190
rect 3012 1180 3078 1190
rect 3204 1180 3270 1190
rect 3688 1180 3754 1190
rect 3880 1180 3946 1190
rect 4072 1180 4138 1190
rect 4264 1180 4330 1190
rect 4456 1180 4522 1190
rect 4648 1180 4714 1190
rect 4840 1180 4906 1190
rect 5032 1180 5098 1190
rect 5516 1180 5582 1190
rect 5708 1180 5774 1190
rect 5900 1180 5966 1190
rect 6092 1180 6158 1190
rect 6284 1180 6350 1190
rect 6476 1180 6542 1190
rect 6668 1180 6734 1190
rect 6860 1180 6926 1190
rect 7344 1180 7410 1190
rect 7536 1180 7602 1190
rect 7728 1180 7794 1190
rect 7920 1180 7986 1190
rect 8112 1180 8178 1190
rect 8304 1180 8370 1190
rect 8496 1180 8562 1190
rect 8688 1180 8754 1190
rect 9172 1180 9238 1190
rect 9364 1180 9430 1190
rect 9556 1180 9622 1190
rect 9748 1180 9814 1190
rect 9940 1180 10006 1190
rect 10132 1180 10198 1190
rect 10324 1180 10390 1190
rect 10516 1180 10582 1190
rect 11000 1180 11066 1190
rect 11192 1180 11258 1190
rect 11384 1180 11450 1190
rect 11576 1180 11642 1190
rect 11768 1180 11834 1190
rect 11960 1180 12026 1190
rect 12152 1180 12218 1190
rect 12344 1180 12410 1190
rect 12828 1180 12894 1190
rect 13020 1180 13086 1190
rect 13212 1180 13278 1190
rect 13404 1180 13470 1190
rect 13596 1180 13662 1190
rect 13788 1180 13854 1190
rect 13980 1180 14046 1190
rect 14172 1180 14238 1190
rect 14656 1180 14722 1190
rect 14848 1180 14914 1190
rect 15040 1180 15106 1190
rect 15232 1180 15298 1190
rect 15424 1180 15490 1190
rect 15616 1180 15682 1190
rect 15808 1180 15874 1190
rect 16000 1180 16066 1190
rect 16484 1180 16550 1190
rect 16676 1180 16742 1190
rect 16868 1180 16934 1190
rect 17060 1180 17126 1190
rect 17252 1180 17318 1190
rect 17444 1180 17510 1190
rect 17636 1180 17702 1190
rect 17828 1180 17894 1190
rect 18312 1180 18378 1190
rect 18504 1180 18570 1190
rect 18696 1180 18762 1190
rect 18888 1180 18954 1190
rect 19080 1180 19146 1190
rect 19272 1180 19338 1190
rect 19464 1180 19530 1190
rect 19656 1180 19722 1190
rect 20140 1180 20206 1190
rect 20332 1180 20398 1190
rect 20524 1180 20590 1190
rect 20716 1180 20782 1190
rect 20908 1180 20974 1190
rect 21100 1180 21166 1190
rect 21292 1180 21358 1190
rect 21484 1180 21550 1190
rect 0 1027 32 1180
rect 98 1027 224 1180
rect 290 1027 416 1180
rect 482 1027 608 1180
rect 674 1027 800 1180
rect 866 1027 992 1180
rect 1058 1027 1184 1180
rect 1250 1027 1376 1180
rect 1828 1027 1860 1180
rect 1926 1027 2052 1180
rect 2118 1027 2244 1180
rect 2310 1027 2436 1180
rect 2502 1027 2628 1180
rect 2694 1027 2820 1180
rect 2886 1027 3012 1180
rect 3078 1027 3204 1180
rect 3656 1027 3688 1180
rect 3754 1027 3880 1180
rect 3946 1027 4072 1180
rect 4138 1027 4264 1180
rect 4330 1027 4456 1180
rect 4522 1027 4648 1180
rect 4714 1027 4840 1180
rect 4906 1027 5032 1180
rect 5484 1027 5516 1180
rect 5582 1027 5708 1180
rect 5774 1027 5900 1180
rect 5966 1027 6092 1180
rect 6158 1027 6284 1180
rect 6350 1027 6476 1180
rect 6542 1027 6668 1180
rect 6734 1027 6860 1180
rect 7312 1027 7344 1180
rect 7410 1027 7536 1180
rect 7602 1027 7728 1180
rect 7794 1027 7920 1180
rect 7986 1027 8112 1180
rect 8178 1027 8304 1180
rect 8370 1027 8496 1180
rect 8562 1027 8688 1180
rect 9140 1027 9172 1180
rect 9238 1027 9364 1180
rect 9430 1027 9556 1180
rect 9622 1027 9748 1180
rect 9814 1027 9940 1180
rect 10006 1027 10132 1180
rect 10198 1027 10324 1180
rect 10390 1027 10516 1180
rect 10968 1027 11000 1180
rect 11066 1027 11192 1180
rect 11258 1027 11384 1180
rect 11450 1027 11576 1180
rect 11642 1027 11768 1180
rect 11834 1027 11960 1180
rect 12026 1027 12152 1180
rect 12218 1027 12344 1180
rect 12796 1027 12828 1180
rect 12894 1027 13020 1180
rect 13086 1027 13212 1180
rect 13278 1027 13404 1180
rect 13470 1027 13596 1180
rect 13662 1027 13788 1180
rect 13854 1027 13980 1180
rect 14046 1027 14172 1180
rect 14624 1027 14656 1180
rect 14722 1027 14848 1180
rect 14914 1027 15040 1180
rect 15106 1027 15232 1180
rect 15298 1027 15424 1180
rect 15490 1027 15616 1180
rect 15682 1027 15808 1180
rect 15874 1027 16000 1180
rect 16452 1027 16484 1180
rect 16550 1027 16676 1180
rect 16742 1027 16868 1180
rect 16934 1027 17060 1180
rect 17126 1027 17252 1180
rect 17318 1027 17444 1180
rect 17510 1027 17636 1180
rect 17702 1027 17828 1180
rect 18280 1027 18312 1180
rect 18378 1027 18504 1180
rect 18570 1027 18696 1180
rect 18762 1027 18888 1180
rect 18954 1027 19080 1180
rect 19146 1027 19272 1180
rect 19338 1027 19464 1180
rect 19530 1027 19656 1180
rect 20108 1027 20140 1180
rect 20206 1027 20332 1180
rect 20398 1027 20524 1180
rect 20590 1027 20716 1180
rect 20782 1027 20908 1180
rect 20974 1027 21100 1180
rect 21166 1027 21292 1180
rect 21358 1027 21484 1180
rect 32 1017 98 1027
rect 224 1017 290 1027
rect 416 1017 482 1027
rect 608 1017 674 1027
rect 800 1017 866 1027
rect 992 1017 1058 1027
rect 1184 1017 1250 1027
rect 1376 1017 1442 1027
rect 1860 1017 1926 1027
rect 2052 1017 2118 1027
rect 2244 1017 2310 1027
rect 2436 1017 2502 1027
rect 2628 1017 2694 1027
rect 2820 1017 2886 1027
rect 3012 1017 3078 1027
rect 3204 1017 3270 1027
rect 3688 1017 3754 1027
rect 3880 1017 3946 1027
rect 4072 1017 4138 1027
rect 4264 1017 4330 1027
rect 4456 1017 4522 1027
rect 4648 1017 4714 1027
rect 4840 1017 4906 1027
rect 5032 1017 5098 1027
rect 5516 1017 5582 1027
rect 5708 1017 5774 1027
rect 5900 1017 5966 1027
rect 6092 1017 6158 1027
rect 6284 1017 6350 1027
rect 6476 1017 6542 1027
rect 6668 1017 6734 1027
rect 6860 1017 6926 1027
rect 7344 1017 7410 1027
rect 7536 1017 7602 1027
rect 7728 1017 7794 1027
rect 7920 1017 7986 1027
rect 8112 1017 8178 1027
rect 8304 1017 8370 1027
rect 8496 1017 8562 1027
rect 8688 1017 8754 1027
rect 9172 1017 9238 1027
rect 9364 1017 9430 1027
rect 9556 1017 9622 1027
rect 9748 1017 9814 1027
rect 9940 1017 10006 1027
rect 10132 1017 10198 1027
rect 10324 1017 10390 1027
rect 10516 1017 10582 1027
rect 11000 1017 11066 1027
rect 11192 1017 11258 1027
rect 11384 1017 11450 1027
rect 11576 1017 11642 1027
rect 11768 1017 11834 1027
rect 11960 1017 12026 1027
rect 12152 1017 12218 1027
rect 12344 1017 12410 1027
rect 12828 1017 12894 1027
rect 13020 1017 13086 1027
rect 13212 1017 13278 1027
rect 13404 1017 13470 1027
rect 13596 1017 13662 1027
rect 13788 1017 13854 1027
rect 13980 1017 14046 1027
rect 14172 1017 14238 1027
rect 14656 1017 14722 1027
rect 14848 1017 14914 1027
rect 15040 1017 15106 1027
rect 15232 1017 15298 1027
rect 15424 1017 15490 1027
rect 15616 1017 15682 1027
rect 15808 1017 15874 1027
rect 16000 1017 16066 1027
rect 16484 1017 16550 1027
rect 16676 1017 16742 1027
rect 16868 1017 16934 1027
rect 17060 1017 17126 1027
rect 17252 1017 17318 1027
rect 17444 1017 17510 1027
rect 17636 1017 17702 1027
rect 17828 1017 17894 1027
rect 18312 1017 18378 1027
rect 18504 1017 18570 1027
rect 18696 1017 18762 1027
rect 18888 1017 18954 1027
rect 19080 1017 19146 1027
rect 19272 1017 19338 1027
rect 19464 1017 19530 1027
rect 19656 1017 19722 1027
rect 20140 1017 20206 1027
rect 20332 1017 20398 1027
rect 20524 1017 20590 1027
rect 20716 1017 20782 1027
rect 20908 1017 20974 1027
rect 21100 1017 21166 1027
rect 21292 1017 21358 1027
rect 21484 1017 21550 1027
rect 128 967 194 977
rect 320 967 386 977
rect 512 967 578 977
rect 704 967 770 977
rect 896 967 962 977
rect 1088 967 1154 977
rect 1280 967 1346 977
rect 1472 967 1528 977
rect 1956 967 2022 977
rect 2148 967 2214 977
rect 2340 967 2406 977
rect 2532 967 2598 977
rect 2724 967 2790 977
rect 2916 967 2982 977
rect 3108 967 3174 977
rect 3300 967 3356 977
rect 3784 967 3850 977
rect 3976 967 4042 977
rect 4168 967 4234 977
rect 4360 967 4426 977
rect 4552 967 4618 977
rect 4744 967 4810 977
rect 4936 967 5002 977
rect 5128 967 5184 977
rect 5612 967 5678 977
rect 5804 967 5870 977
rect 5996 967 6062 977
rect 6188 967 6254 977
rect 6380 967 6446 977
rect 6572 967 6638 977
rect 6764 967 6830 977
rect 6956 967 7012 977
rect 7440 967 7506 977
rect 7632 967 7698 977
rect 7824 967 7890 977
rect 8016 967 8082 977
rect 8208 967 8274 977
rect 8400 967 8466 977
rect 8592 967 8658 977
rect 8784 967 8840 977
rect 9268 967 9334 977
rect 9460 967 9526 977
rect 9652 967 9718 977
rect 9844 967 9910 977
rect 10036 967 10102 977
rect 10228 967 10294 977
rect 10420 967 10486 977
rect 10612 967 10668 977
rect 11096 967 11162 977
rect 11288 967 11354 977
rect 11480 967 11546 977
rect 11672 967 11738 977
rect 11864 967 11930 977
rect 12056 967 12122 977
rect 12248 967 12314 977
rect 12440 967 12496 977
rect 12924 967 12990 977
rect 13116 967 13182 977
rect 13308 967 13374 977
rect 13500 967 13566 977
rect 13692 967 13758 977
rect 13884 967 13950 977
rect 14076 967 14142 977
rect 14268 967 14324 977
rect 14752 967 14818 977
rect 14944 967 15010 977
rect 15136 967 15202 977
rect 15328 967 15394 977
rect 15520 967 15586 977
rect 15712 967 15778 977
rect 15904 967 15970 977
rect 16096 967 16152 977
rect 16580 967 16646 977
rect 16772 967 16838 977
rect 16964 967 17030 977
rect 17156 967 17222 977
rect 17348 967 17414 977
rect 17540 967 17606 977
rect 17732 967 17798 977
rect 17924 967 17980 977
rect 18408 967 18474 977
rect 18600 967 18666 977
rect 18792 967 18858 977
rect 18984 967 19050 977
rect 19176 967 19242 977
rect 19368 967 19434 977
rect 19560 967 19626 977
rect 19752 967 19808 977
rect 20236 967 20302 977
rect 20428 967 20494 977
rect 20620 967 20686 977
rect 20812 967 20878 977
rect 21004 967 21070 977
rect 21196 967 21262 977
rect 21388 967 21454 977
rect 21580 967 21636 977
rect 0 814 128 967
rect 194 814 320 967
rect 386 814 512 967
rect 578 814 704 967
rect 770 814 896 967
rect 962 814 1088 967
rect 1154 814 1280 967
rect 1346 814 1472 967
rect 1528 814 1708 967
rect 1828 814 1956 967
rect 2022 814 2148 967
rect 2214 814 2340 967
rect 2406 814 2532 967
rect 2598 814 2724 967
rect 2790 814 2916 967
rect 2982 814 3108 967
rect 3174 814 3300 967
rect 3356 814 3536 967
rect 3656 814 3784 967
rect 3850 814 3976 967
rect 4042 814 4168 967
rect 4234 814 4360 967
rect 4426 814 4552 967
rect 4618 814 4744 967
rect 4810 814 4936 967
rect 5002 814 5128 967
rect 5184 814 5364 967
rect 5484 814 5612 967
rect 5678 814 5804 967
rect 5870 814 5996 967
rect 6062 814 6188 967
rect 6254 814 6380 967
rect 6446 814 6572 967
rect 6638 814 6764 967
rect 6830 814 6956 967
rect 7012 814 7192 967
rect 7312 814 7440 967
rect 7506 814 7632 967
rect 7698 814 7824 967
rect 7890 814 8016 967
rect 8082 814 8208 967
rect 8274 814 8400 967
rect 8466 814 8592 967
rect 8658 814 8784 967
rect 8840 814 9020 967
rect 9140 814 9268 967
rect 9334 814 9460 967
rect 9526 814 9652 967
rect 9718 814 9844 967
rect 9910 814 10036 967
rect 10102 814 10228 967
rect 10294 814 10420 967
rect 10486 814 10612 967
rect 10668 814 10848 967
rect 10968 814 11096 967
rect 11162 814 11288 967
rect 11354 814 11480 967
rect 11546 814 11672 967
rect 11738 814 11864 967
rect 11930 814 12056 967
rect 12122 814 12248 967
rect 12314 814 12440 967
rect 12496 814 12676 967
rect 12796 814 12924 967
rect 12990 814 13116 967
rect 13182 814 13308 967
rect 13374 814 13500 967
rect 13566 814 13692 967
rect 13758 814 13884 967
rect 13950 814 14076 967
rect 14142 814 14268 967
rect 14324 814 14504 967
rect 14624 814 14752 967
rect 14818 814 14944 967
rect 15010 814 15136 967
rect 15202 814 15328 967
rect 15394 814 15520 967
rect 15586 814 15712 967
rect 15778 814 15904 967
rect 15970 814 16096 967
rect 16152 814 16332 967
rect 16452 814 16580 967
rect 16646 814 16772 967
rect 16838 814 16964 967
rect 17030 814 17156 967
rect 17222 814 17348 967
rect 17414 814 17540 967
rect 17606 814 17732 967
rect 17798 814 17924 967
rect 17980 814 18160 967
rect 18280 814 18408 967
rect 18474 814 18600 967
rect 18666 814 18792 967
rect 18858 814 18984 967
rect 19050 814 19176 967
rect 19242 814 19368 967
rect 19434 814 19560 967
rect 19626 814 19752 967
rect 19808 814 19988 967
rect 20108 814 20236 967
rect 20302 814 20428 967
rect 20494 814 20620 967
rect 20686 814 20812 967
rect 20878 814 21004 967
rect 21070 814 21196 967
rect 21262 814 21388 967
rect 21454 814 21580 967
rect 21636 814 21816 967
rect 128 804 194 814
rect 320 804 386 814
rect 512 804 578 814
rect 704 804 770 814
rect 896 804 962 814
rect 1088 804 1154 814
rect 1280 804 1346 814
rect 1472 804 1528 814
rect 1956 804 2022 814
rect 2148 804 2214 814
rect 2340 804 2406 814
rect 2532 804 2598 814
rect 2724 804 2790 814
rect 2916 804 2982 814
rect 3108 804 3174 814
rect 3300 804 3356 814
rect 3784 804 3850 814
rect 3976 804 4042 814
rect 4168 804 4234 814
rect 4360 804 4426 814
rect 4552 804 4618 814
rect 4744 804 4810 814
rect 4936 804 5002 814
rect 5128 804 5184 814
rect 5612 804 5678 814
rect 5804 804 5870 814
rect 5996 804 6062 814
rect 6188 804 6254 814
rect 6380 804 6446 814
rect 6572 804 6638 814
rect 6764 804 6830 814
rect 6956 804 7012 814
rect 7440 804 7506 814
rect 7632 804 7698 814
rect 7824 804 7890 814
rect 8016 804 8082 814
rect 8208 804 8274 814
rect 8400 804 8466 814
rect 8592 804 8658 814
rect 8784 804 8840 814
rect 9268 804 9334 814
rect 9460 804 9526 814
rect 9652 804 9718 814
rect 9844 804 9910 814
rect 10036 804 10102 814
rect 10228 804 10294 814
rect 10420 804 10486 814
rect 10612 804 10668 814
rect 11096 804 11162 814
rect 11288 804 11354 814
rect 11480 804 11546 814
rect 11672 804 11738 814
rect 11864 804 11930 814
rect 12056 804 12122 814
rect 12248 804 12314 814
rect 12440 804 12496 814
rect 12924 804 12990 814
rect 13116 804 13182 814
rect 13308 804 13374 814
rect 13500 804 13566 814
rect 13692 804 13758 814
rect 13884 804 13950 814
rect 14076 804 14142 814
rect 14268 804 14324 814
rect 14752 804 14818 814
rect 14944 804 15010 814
rect 15136 804 15202 814
rect 15328 804 15394 814
rect 15520 804 15586 814
rect 15712 804 15778 814
rect 15904 804 15970 814
rect 16096 804 16152 814
rect 16580 804 16646 814
rect 16772 804 16838 814
rect 16964 804 17030 814
rect 17156 804 17222 814
rect 17348 804 17414 814
rect 17540 804 17606 814
rect 17732 804 17798 814
rect 17924 804 17980 814
rect 18408 804 18474 814
rect 18600 804 18666 814
rect 18792 804 18858 814
rect 18984 804 19050 814
rect 19176 804 19242 814
rect 19368 804 19434 814
rect 19560 804 19626 814
rect 19752 804 19808 814
rect 20236 804 20302 814
rect 20428 804 20494 814
rect 20620 804 20686 814
rect 20812 804 20878 814
rect 21004 804 21070 814
rect 21196 804 21262 814
rect 21388 804 21454 814
rect 21580 804 21636 814
rect 32 466 98 476
rect 224 466 290 476
rect 416 466 482 476
rect 608 466 674 476
rect 800 466 866 476
rect 992 466 1058 476
rect 1184 466 1250 476
rect 1376 466 1442 476
rect 1860 466 1926 476
rect 2052 466 2118 476
rect 2244 466 2310 476
rect 2436 466 2502 476
rect 2628 466 2694 476
rect 2820 466 2886 476
rect 3012 466 3078 476
rect 3204 466 3270 476
rect 3688 466 3754 476
rect 3880 466 3946 476
rect 4072 466 4138 476
rect 4264 466 4330 476
rect 4456 466 4522 476
rect 4648 466 4714 476
rect 4840 466 4906 476
rect 5032 466 5098 476
rect 5516 466 5582 476
rect 5708 466 5774 476
rect 5900 466 5966 476
rect 6092 466 6158 476
rect 6284 466 6350 476
rect 6476 466 6542 476
rect 6668 466 6734 476
rect 6860 466 6926 476
rect 7344 466 7410 476
rect 7536 466 7602 476
rect 7728 466 7794 476
rect 7920 466 7986 476
rect 8112 466 8178 476
rect 8304 466 8370 476
rect 8496 466 8562 476
rect 8688 466 8754 476
rect 9172 466 9238 476
rect 9364 466 9430 476
rect 9556 466 9622 476
rect 9748 466 9814 476
rect 9940 466 10006 476
rect 10132 466 10198 476
rect 10324 466 10390 476
rect 10516 466 10582 476
rect 11000 466 11066 476
rect 11192 466 11258 476
rect 11384 466 11450 476
rect 11576 466 11642 476
rect 11768 466 11834 476
rect 11960 466 12026 476
rect 12152 466 12218 476
rect 12344 466 12410 476
rect 12828 466 12894 476
rect 13020 466 13086 476
rect 13212 466 13278 476
rect 13404 466 13470 476
rect 13596 466 13662 476
rect 13788 466 13854 476
rect 13980 466 14046 476
rect 14172 466 14238 476
rect 14656 466 14722 476
rect 14848 466 14914 476
rect 15040 466 15106 476
rect 15232 466 15298 476
rect 15424 466 15490 476
rect 15616 466 15682 476
rect 15808 466 15874 476
rect 16000 466 16066 476
rect 16484 466 16550 476
rect 16676 466 16742 476
rect 16868 466 16934 476
rect 17060 466 17126 476
rect 17252 466 17318 476
rect 17444 466 17510 476
rect 17636 466 17702 476
rect 17828 466 17894 476
rect 18312 466 18378 476
rect 18504 466 18570 476
rect 18696 466 18762 476
rect 18888 466 18954 476
rect 19080 466 19146 476
rect 19272 466 19338 476
rect 19464 466 19530 476
rect 19656 466 19722 476
rect 20140 466 20206 476
rect 20332 466 20398 476
rect 20524 466 20590 476
rect 20716 466 20782 476
rect 20908 466 20974 476
rect 21100 466 21166 476
rect 21292 466 21358 476
rect 21484 466 21550 476
rect 0 313 32 466
rect 98 313 224 466
rect 290 313 416 466
rect 482 313 608 466
rect 674 313 800 466
rect 866 313 992 466
rect 1058 313 1184 466
rect 1250 313 1376 466
rect 1828 313 1860 466
rect 1926 313 2052 466
rect 2118 313 2244 466
rect 2310 313 2436 466
rect 2502 313 2628 466
rect 2694 313 2820 466
rect 2886 313 3012 466
rect 3078 313 3204 466
rect 3656 313 3688 466
rect 3754 313 3880 466
rect 3946 313 4072 466
rect 4138 313 4264 466
rect 4330 313 4456 466
rect 4522 313 4648 466
rect 4714 313 4840 466
rect 4906 313 5032 466
rect 5484 313 5516 466
rect 5582 313 5708 466
rect 5774 313 5900 466
rect 5966 313 6092 466
rect 6158 313 6284 466
rect 6350 313 6476 466
rect 6542 313 6668 466
rect 6734 313 6860 466
rect 7312 313 7344 466
rect 7410 313 7536 466
rect 7602 313 7728 466
rect 7794 313 7920 466
rect 7986 313 8112 466
rect 8178 313 8304 466
rect 8370 313 8496 466
rect 8562 313 8688 466
rect 9140 313 9172 466
rect 9238 313 9364 466
rect 9430 313 9556 466
rect 9622 313 9748 466
rect 9814 313 9940 466
rect 10006 313 10132 466
rect 10198 313 10324 466
rect 10390 313 10516 466
rect 10968 313 11000 466
rect 11066 313 11192 466
rect 11258 313 11384 466
rect 11450 313 11576 466
rect 11642 313 11768 466
rect 11834 313 11960 466
rect 12026 313 12152 466
rect 12218 313 12344 466
rect 12796 313 12828 466
rect 12894 313 13020 466
rect 13086 313 13212 466
rect 13278 313 13404 466
rect 13470 313 13596 466
rect 13662 313 13788 466
rect 13854 313 13980 466
rect 14046 313 14172 466
rect 14624 313 14656 466
rect 14722 313 14848 466
rect 14914 313 15040 466
rect 15106 313 15232 466
rect 15298 313 15424 466
rect 15490 313 15616 466
rect 15682 313 15808 466
rect 15874 313 16000 466
rect 16452 313 16484 466
rect 16550 313 16676 466
rect 16742 313 16868 466
rect 16934 313 17060 466
rect 17126 313 17252 466
rect 17318 313 17444 466
rect 17510 313 17636 466
rect 17702 313 17828 466
rect 18280 313 18312 466
rect 18378 313 18504 466
rect 18570 313 18696 466
rect 18762 313 18888 466
rect 18954 313 19080 466
rect 19146 313 19272 466
rect 19338 313 19464 466
rect 19530 313 19656 466
rect 20108 313 20140 466
rect 20206 313 20332 466
rect 20398 313 20524 466
rect 20590 313 20716 466
rect 20782 313 20908 466
rect 20974 313 21100 466
rect 21166 313 21292 466
rect 21358 313 21484 466
rect 32 303 98 313
rect 224 303 290 313
rect 416 303 482 313
rect 608 303 674 313
rect 800 303 866 313
rect 992 303 1058 313
rect 1184 303 1250 313
rect 1376 303 1442 313
rect 1860 303 1926 313
rect 2052 303 2118 313
rect 2244 303 2310 313
rect 2436 303 2502 313
rect 2628 303 2694 313
rect 2820 303 2886 313
rect 3012 303 3078 313
rect 3204 303 3270 313
rect 3688 303 3754 313
rect 3880 303 3946 313
rect 4072 303 4138 313
rect 4264 303 4330 313
rect 4456 303 4522 313
rect 4648 303 4714 313
rect 4840 303 4906 313
rect 5032 303 5098 313
rect 5516 303 5582 313
rect 5708 303 5774 313
rect 5900 303 5966 313
rect 6092 303 6158 313
rect 6284 303 6350 313
rect 6476 303 6542 313
rect 6668 303 6734 313
rect 6860 303 6926 313
rect 7344 303 7410 313
rect 7536 303 7602 313
rect 7728 303 7794 313
rect 7920 303 7986 313
rect 8112 303 8178 313
rect 8304 303 8370 313
rect 8496 303 8562 313
rect 8688 303 8754 313
rect 9172 303 9238 313
rect 9364 303 9430 313
rect 9556 303 9622 313
rect 9748 303 9814 313
rect 9940 303 10006 313
rect 10132 303 10198 313
rect 10324 303 10390 313
rect 10516 303 10582 313
rect 11000 303 11066 313
rect 11192 303 11258 313
rect 11384 303 11450 313
rect 11576 303 11642 313
rect 11768 303 11834 313
rect 11960 303 12026 313
rect 12152 303 12218 313
rect 12344 303 12410 313
rect 12828 303 12894 313
rect 13020 303 13086 313
rect 13212 303 13278 313
rect 13404 303 13470 313
rect 13596 303 13662 313
rect 13788 303 13854 313
rect 13980 303 14046 313
rect 14172 303 14238 313
rect 14656 303 14722 313
rect 14848 303 14914 313
rect 15040 303 15106 313
rect 15232 303 15298 313
rect 15424 303 15490 313
rect 15616 303 15682 313
rect 15808 303 15874 313
rect 16000 303 16066 313
rect 16484 303 16550 313
rect 16676 303 16742 313
rect 16868 303 16934 313
rect 17060 303 17126 313
rect 17252 303 17318 313
rect 17444 303 17510 313
rect 17636 303 17702 313
rect 17828 303 17894 313
rect 18312 303 18378 313
rect 18504 303 18570 313
rect 18696 303 18762 313
rect 18888 303 18954 313
rect 19080 303 19146 313
rect 19272 303 19338 313
rect 19464 303 19530 313
rect 19656 303 19722 313
rect 20140 303 20206 313
rect 20332 303 20398 313
rect 20524 303 20590 313
rect 20716 303 20782 313
rect 20908 303 20974 313
rect 21100 303 21166 313
rect 21292 303 21358 313
rect 21484 303 21550 313
rect 128 253 194 263
rect 320 253 386 263
rect 512 253 578 263
rect 704 253 770 263
rect 896 253 962 263
rect 1088 253 1154 263
rect 1280 253 1346 263
rect 1472 253 1528 263
rect 1956 253 2022 263
rect 2148 253 2214 263
rect 2340 253 2406 263
rect 2532 253 2598 263
rect 2724 253 2790 263
rect 2916 253 2982 263
rect 3108 253 3174 263
rect 3300 253 3356 263
rect 3784 253 3850 263
rect 3976 253 4042 263
rect 4168 253 4234 263
rect 4360 253 4426 263
rect 4552 253 4618 263
rect 4744 253 4810 263
rect 4936 253 5002 263
rect 5128 253 5184 263
rect 5612 253 5678 263
rect 5804 253 5870 263
rect 5996 253 6062 263
rect 6188 253 6254 263
rect 6380 253 6446 263
rect 6572 253 6638 263
rect 6764 253 6830 263
rect 6956 253 7012 263
rect 7440 253 7506 263
rect 7632 253 7698 263
rect 7824 253 7890 263
rect 8016 253 8082 263
rect 8208 253 8274 263
rect 8400 253 8466 263
rect 8592 253 8658 263
rect 8784 253 8840 263
rect 9268 253 9334 263
rect 9460 253 9526 263
rect 9652 253 9718 263
rect 9844 253 9910 263
rect 10036 253 10102 263
rect 10228 253 10294 263
rect 10420 253 10486 263
rect 10612 253 10668 263
rect 11096 253 11162 263
rect 11288 253 11354 263
rect 11480 253 11546 263
rect 11672 253 11738 263
rect 11864 253 11930 263
rect 12056 253 12122 263
rect 12248 253 12314 263
rect 12440 253 12496 263
rect 12924 253 12990 263
rect 13116 253 13182 263
rect 13308 253 13374 263
rect 13500 253 13566 263
rect 13692 253 13758 263
rect 13884 253 13950 263
rect 14076 253 14142 263
rect 14268 253 14324 263
rect 14752 253 14818 263
rect 14944 253 15010 263
rect 15136 253 15202 263
rect 15328 253 15394 263
rect 15520 253 15586 263
rect 15712 253 15778 263
rect 15904 253 15970 263
rect 16096 253 16152 263
rect 16580 253 16646 263
rect 16772 253 16838 263
rect 16964 253 17030 263
rect 17156 253 17222 263
rect 17348 253 17414 263
rect 17540 253 17606 263
rect 17732 253 17798 263
rect 17924 253 17980 263
rect 18408 253 18474 263
rect 18600 253 18666 263
rect 18792 253 18858 263
rect 18984 253 19050 263
rect 19176 253 19242 263
rect 19368 253 19434 263
rect 19560 253 19626 263
rect 19752 253 19808 263
rect 20236 253 20302 263
rect 20428 253 20494 263
rect 20620 253 20686 263
rect 20812 253 20878 263
rect 21004 253 21070 263
rect 21196 253 21262 263
rect 21388 253 21454 263
rect 21580 253 21636 263
rect 0 100 128 253
rect 194 100 320 253
rect 386 100 512 253
rect 578 100 704 253
rect 770 100 896 253
rect 962 100 1088 253
rect 1154 100 1280 253
rect 1346 100 1472 253
rect 1528 100 1708 253
rect 1828 100 1956 253
rect 2022 100 2148 253
rect 2214 100 2340 253
rect 2406 100 2532 253
rect 2598 100 2724 253
rect 2790 100 2916 253
rect 2982 100 3108 253
rect 3174 100 3300 253
rect 3356 100 3536 253
rect 3656 100 3784 253
rect 3850 100 3976 253
rect 4042 100 4168 253
rect 4234 100 4360 253
rect 4426 100 4552 253
rect 4618 100 4744 253
rect 4810 100 4936 253
rect 5002 100 5128 253
rect 5184 100 5364 253
rect 5484 100 5612 253
rect 5678 100 5804 253
rect 5870 100 5996 253
rect 6062 100 6188 253
rect 6254 100 6380 253
rect 6446 100 6572 253
rect 6638 100 6764 253
rect 6830 100 6956 253
rect 7012 100 7192 253
rect 7312 100 7440 253
rect 7506 100 7632 253
rect 7698 100 7824 253
rect 7890 100 8016 253
rect 8082 100 8208 253
rect 8274 100 8400 253
rect 8466 100 8592 253
rect 8658 100 8784 253
rect 8840 100 9020 253
rect 9140 100 9268 253
rect 9334 100 9460 253
rect 9526 100 9652 253
rect 9718 100 9844 253
rect 9910 100 10036 253
rect 10102 100 10228 253
rect 10294 100 10420 253
rect 10486 100 10612 253
rect 10668 100 10848 253
rect 10968 100 11096 253
rect 11162 100 11288 253
rect 11354 100 11480 253
rect 11546 100 11672 253
rect 11738 100 11864 253
rect 11930 100 12056 253
rect 12122 100 12248 253
rect 12314 100 12440 253
rect 12496 100 12676 253
rect 12796 100 12924 253
rect 12990 100 13116 253
rect 13182 100 13308 253
rect 13374 100 13500 253
rect 13566 100 13692 253
rect 13758 100 13884 253
rect 13950 100 14076 253
rect 14142 100 14268 253
rect 14324 100 14504 253
rect 14624 100 14752 253
rect 14818 100 14944 253
rect 15010 100 15136 253
rect 15202 100 15328 253
rect 15394 100 15520 253
rect 15586 100 15712 253
rect 15778 100 15904 253
rect 15970 100 16096 253
rect 16152 100 16332 253
rect 16452 100 16580 253
rect 16646 100 16772 253
rect 16838 100 16964 253
rect 17030 100 17156 253
rect 17222 100 17348 253
rect 17414 100 17540 253
rect 17606 100 17732 253
rect 17798 100 17924 253
rect 17980 100 18160 253
rect 18280 100 18408 253
rect 18474 100 18600 253
rect 18666 100 18792 253
rect 18858 100 18984 253
rect 19050 100 19176 253
rect 19242 100 19368 253
rect 19434 100 19560 253
rect 19626 100 19752 253
rect 19808 100 19988 253
rect 20108 100 20236 253
rect 20302 100 20428 253
rect 20494 100 20620 253
rect 20686 100 20812 253
rect 20878 100 21004 253
rect 21070 100 21196 253
rect 21262 100 21388 253
rect 21454 100 21580 253
rect 21636 100 21816 253
rect 128 90 194 100
rect 320 90 386 100
rect 512 90 578 100
rect 704 90 770 100
rect 896 90 962 100
rect 1088 90 1154 100
rect 1280 90 1346 100
rect 1472 90 1528 100
rect 1956 90 2022 100
rect 2148 90 2214 100
rect 2340 90 2406 100
rect 2532 90 2598 100
rect 2724 90 2790 100
rect 2916 90 2982 100
rect 3108 90 3174 100
rect 3300 90 3356 100
rect 3784 90 3850 100
rect 3976 90 4042 100
rect 4168 90 4234 100
rect 4360 90 4426 100
rect 4552 90 4618 100
rect 4744 90 4810 100
rect 4936 90 5002 100
rect 5128 90 5184 100
rect 5612 90 5678 100
rect 5804 90 5870 100
rect 5996 90 6062 100
rect 6188 90 6254 100
rect 6380 90 6446 100
rect 6572 90 6638 100
rect 6764 90 6830 100
rect 6956 90 7012 100
rect 7440 90 7506 100
rect 7632 90 7698 100
rect 7824 90 7890 100
rect 8016 90 8082 100
rect 8208 90 8274 100
rect 8400 90 8466 100
rect 8592 90 8658 100
rect 8784 90 8840 100
rect 9268 90 9334 100
rect 9460 90 9526 100
rect 9652 90 9718 100
rect 9844 90 9910 100
rect 10036 90 10102 100
rect 10228 90 10294 100
rect 10420 90 10486 100
rect 10612 90 10668 100
rect 11096 90 11162 100
rect 11288 90 11354 100
rect 11480 90 11546 100
rect 11672 90 11738 100
rect 11864 90 11930 100
rect 12056 90 12122 100
rect 12248 90 12314 100
rect 12440 90 12496 100
rect 12924 90 12990 100
rect 13116 90 13182 100
rect 13308 90 13374 100
rect 13500 90 13566 100
rect 13692 90 13758 100
rect 13884 90 13950 100
rect 14076 90 14142 100
rect 14268 90 14324 100
rect 14752 90 14818 100
rect 14944 90 15010 100
rect 15136 90 15202 100
rect 15328 90 15394 100
rect 15520 90 15586 100
rect 15712 90 15778 100
rect 15904 90 15970 100
rect 16096 90 16152 100
rect 16580 90 16646 100
rect 16772 90 16838 100
rect 16964 90 17030 100
rect 17156 90 17222 100
rect 17348 90 17414 100
rect 17540 90 17606 100
rect 17732 90 17798 100
rect 17924 90 17980 100
rect 18408 90 18474 100
rect 18600 90 18666 100
rect 18792 90 18858 100
rect 18984 90 19050 100
rect 19176 90 19242 100
rect 19368 90 19434 100
rect 19560 90 19626 100
rect 19752 90 19808 100
rect 20236 90 20302 100
rect 20428 90 20494 100
rect 20620 90 20686 100
rect 20812 90 20878 100
rect 21004 90 21070 100
rect 21196 90 21262 100
rect 21388 90 21454 100
rect 21580 90 21636 100
use sky130_fd_pr__pfet_01v8_KPD88M  sky130_fd_pr__pfet_01v8_KPD88M_0
array 0 11 1828 0 29 714
timestamp 1697921066
transform 1 0 785 0 1 300
box -785 -300 785 300
<< end >>
