magic
tech sky130A
magscale 1 2
timestamp 1697794388
<< nwell >>
rect -655 -462 655 462
<< pmos >>
rect -561 -400 -501 400
rect -443 -400 -383 400
rect -325 -400 -265 400
rect -207 -400 -147 400
rect -89 -400 -29 400
rect 29 -400 89 400
rect 147 -400 207 400
rect 265 -400 325 400
rect 383 -400 443 400
rect 501 -400 561 400
<< pdiff >>
rect -619 388 -561 400
rect -619 -388 -607 388
rect -573 -388 -561 388
rect -619 -400 -561 -388
rect -501 388 -443 400
rect -501 -388 -489 388
rect -455 -388 -443 388
rect -501 -400 -443 -388
rect -383 388 -325 400
rect -383 -388 -371 388
rect -337 -388 -325 388
rect -383 -400 -325 -388
rect -265 388 -207 400
rect -265 -388 -253 388
rect -219 -388 -207 388
rect -265 -400 -207 -388
rect -147 388 -89 400
rect -147 -388 -135 388
rect -101 -388 -89 388
rect -147 -400 -89 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 89 388 147 400
rect 89 -388 101 388
rect 135 -388 147 388
rect 89 -400 147 -388
rect 207 388 265 400
rect 207 -388 219 388
rect 253 -388 265 388
rect 207 -400 265 -388
rect 325 388 383 400
rect 325 -388 337 388
rect 371 -388 383 388
rect 325 -400 383 -388
rect 443 388 501 400
rect 443 -388 455 388
rect 489 -388 501 388
rect 443 -400 501 -388
rect 561 388 619 400
rect 561 -388 573 388
rect 607 -388 619 388
rect 561 -400 619 -388
<< pdiffc >>
rect -607 -388 -573 388
rect -489 -388 -455 388
rect -371 -388 -337 388
rect -253 -388 -219 388
rect -135 -388 -101 388
rect -17 -388 17 388
rect 101 -388 135 388
rect 219 -388 253 388
rect 337 -388 371 388
rect 455 -388 489 388
rect 573 -388 607 388
<< poly >>
rect -561 400 -501 426
rect -443 400 -383 426
rect -325 400 -265 426
rect -207 400 -147 426
rect -89 400 -29 426
rect 29 400 89 426
rect 147 400 207 426
rect 265 400 325 426
rect 383 400 443 426
rect 501 400 561 426
rect -561 -426 -501 -400
rect -443 -426 -383 -400
rect -325 -426 -265 -400
rect -207 -426 -147 -400
rect -89 -426 -29 -400
rect 29 -426 89 -400
rect 147 -426 207 -400
rect 265 -426 325 -400
rect 383 -426 443 -400
rect 501 -426 561 -400
<< locali >>
rect -607 388 -573 404
rect -607 -404 -573 -388
rect -489 388 -455 404
rect -489 -404 -455 -388
rect -371 388 -337 404
rect -371 -404 -337 -388
rect -253 388 -219 404
rect -253 -404 -219 -388
rect -135 388 -101 404
rect -135 -404 -101 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 101 388 135 404
rect 101 -404 135 -388
rect 219 388 253 404
rect 219 -404 253 -388
rect 337 388 371 404
rect 337 -404 371 -388
rect 455 388 489 404
rect 455 -404 489 -388
rect 573 388 607 404
rect 573 -404 607 -388
<< viali >>
rect -607 -388 -573 388
rect -489 -388 -455 388
rect -371 -388 -337 388
rect -253 -388 -219 388
rect -135 -388 -101 388
rect -17 -388 17 388
rect 101 -388 135 388
rect 219 -388 253 388
rect 337 -388 371 388
rect 455 -388 489 388
rect 573 -388 607 388
<< metal1 >>
rect -613 388 -567 400
rect -613 -388 -607 388
rect -573 -388 -567 388
rect -613 -400 -567 -388
rect -495 388 -449 400
rect -495 -388 -489 388
rect -455 -388 -449 388
rect -495 -400 -449 -388
rect -377 388 -331 400
rect -377 -388 -371 388
rect -337 -388 -331 388
rect -377 -400 -331 -388
rect -259 388 -213 400
rect -259 -388 -253 388
rect -219 -388 -213 388
rect -259 -400 -213 -388
rect -141 388 -95 400
rect -141 -388 -135 388
rect -101 -388 -95 388
rect -141 -400 -95 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 95 388 141 400
rect 95 -388 101 388
rect 135 -388 141 388
rect 95 -400 141 -388
rect 213 388 259 400
rect 213 -388 219 388
rect 253 -388 259 388
rect 213 -400 259 -388
rect 331 388 377 400
rect 331 -388 337 388
rect 371 -388 377 388
rect 331 -400 377 -388
rect 449 388 495 400
rect 449 -388 455 388
rect 489 -388 495 388
rect 449 -400 495 -388
rect 567 388 613 400
rect 567 -388 573 388
rect 607 -388 613 388
rect 567 -400 613 -388
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4 l 0.3 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
